----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:31:20 11/29/2019 
-- Design Name: 
-- Module Name:    ROM_lett_num - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ROM_lett_num is
	Port ( clock, read_enable : in  STD_LOGIC;
           address_x: in  STD_LOGIC_VECTOR (5 downto 0);
			  address_y: in  STD_LOGIC_VECTOR (4 downto 0);
           data_out : out  STD_LOGIC_VECTOR (0 to 31));
end ROM_lett_num;

architecture Behavioral of ROM_lett_num is

type ROM_type is array(0 to 2047) of std_logic_vector(0 to 31);
constant rom : ROM_type := (
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111111111111111111100000",
"00011111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111110000",
"00011111111111111111111111110000",
"00001111111111111111111111000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111111111111111111100000",
"00011111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111111111111111111000000",
"00111111111111111111111111000000",
"00111111111111111111111111000000",
"00111111111111111111111111000000",
"00111111111111111111111111000000",
"00111111111111111111111111000000",
"00111111111111111111111111000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111110000",
"00011111111111111111111111110000",
"00001111111111111111111111000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111000000000111111000000",
"00011111111000000000111111110000",
"00111111111100000000111111110000",
"00111111111100000000111111111000",
"00111111111100000000111111111000",
"00111111111110000000111111111000",
"00111111111110000000111111111000",
"00111111111110000000111111111000",
"00111111111111000000111111111000",
"00111111111111000000111111111000",
"00111111111111000000111111111000",
"00111111111111100000111111111000",
"00111111111111100000111111111000",
"00111111111111100000111111111000",
"00111111111111110000111111111000",
"00111111111111110000111111111000",
"00111111111111110000111111111000",
"00111111111111111000111111111000",
"00111111111111111000111111111000",
"00111111111111111000111111111000",
"00111111111111111100111111111000",
"00111111111111111100111111111000",
"00111111111111111100111111111000",
"00111111111111111110111111111000",
"00111111111111111110111111111000",
"00111111111111111110111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111011111111111111111000",
"00111111111011111111111111111000",
"00111111111011111111111111111000",
"00111111111001111111111111111000",
"00111111111001111111111111111000",
"00111111111000111111111111111000",
"00111111111000111111111111111000",
"00111111111000111111111111111000",
"00111111111000011111111111111000",
"00111111111000011111111111111000",
"00111111111000011111111111111000",
"00111111111000001111111111111000",
"00111111111000001111111111111000",
"00111111111000000111111111111000",
"00111111111000000111111111111000",
"00111111111000000111111111111000",
"00111111111000000011111111111000",
"00111111111000000011111111111000",
"00111111111000000011111111111000",
"00111111111000000001111111111000",
"00111111111000000001111111111000",
"00111111111000000000111111111000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111111111111111111100000",
"00111111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111110000",
"00111111111111111111111111100000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111111111111111111000000",
"00111111111111111111111111100000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111100000",
"00111111111111111111111111000000",
"00111111111000111111110000000000",
"00111111111000111111110000000000",
"00111111111000111111111000000000",
"00111111111000011111111000000000",
"00111111111000011111111000000000",
"00111111111000011111111100000000",
"00111111111000001111111100000000",
"00111111111000001111111110000000",
"00111111111000000111111110000000",
"00111111111000000111111110000000",
"00111111111000000111111111000000",
"00111111111000000011111111000000",
"00111111111000000011111111100000",
"00111111111000000011111111100000",
"00111111111000000001111111110000",
"00111111111000000001111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000011111111100",
"00111111111000000000011111111100",
"00111111111000000000011111111110",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111110000000111111111000",
"00011111111111000000111111111000",
"00011111111111000000111111111000",
"00001111111111000000111111111000",
"00001111111111100000111111111000",
"00000111111111100000111111111000",
"00000111111111110000111111111000",
"00000011111111110000111111111000",
"00000011111111111000111111111000",
"00000011111111111000000000000000",
"00000001111111111100000000000000",
"00000001111111111100000000000000",
"00000000111111111110000000000000",
"00000000111111111110000000000000",
"00000000011111111111000000000000",
"00000000011111111111000000000000",
"00000000001111111111000000000000",
"00000000001111111111100000000000",
"00000000000111111111100000000000",
"00000000000111111111110000000000",
"00000000000011111111110000000000",
"00000000000011111111111000000000",
"00000000000001111111111000000000",
"00000000000001111111111100000000",
"00000000000000111111111100000000",
"00000000000000111111111110000000",
"00111111111000011111111110000000",
"00111111111000011111111110000000",
"00111111111000011111111111000000",
"00111111111000001111111111000000",
"00111111111000001111111111100000",
"00111111111000000111111111100000",
"00111111111000000111111111110000",
"00111111111000000011111111110000",
"00111111111000000011111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111111111111111111111110",
"00111111111111111111111111111110",
"00111111111111111111111111111110",
"00111111111111111111111111111110",
"00111111111111111111111111111110",
"00111111111111111111111111111110",
"00111111111111111111111111111110",
"00111111111111111111111111111110",
"00111111111111111111111111111110",
"00111111111000011111111100000000",
"00111111111000011111111100000000",
"00111111111000011111111100000000",
"00111111111000011111111100000000",
"00111111111000011111111100000000",
"00111111111000011111111100000000",
"00111111111000011111111100000000",
"00111111111000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111000000000111111110000",
"00111111111000000001111111110000",
"00111111111000000001111111110000",
"00111111111000000001111111110000",
"00011111111000000001111111110000",
"00011111111000000001111111110000",
"00011111111100000001111111100000",
"00011111111100000001111111100000",
"00011111111100000001111111100000",
"00011111111100000011111111100000",
"00001111111100000011111111100000",
"00001111111100000011111111100000",
"00001111111100000011111111000000",
"00001111111100000011111111000000",
"00001111111110000011111111000000",
"00001111111110000011111111000000",
"00000111111110000011111111000000",
"00000111111110000111111111000000",
"00000111111110000111111110000000",
"00000111111110000111111110000000",
"00000111111110000111111110000000",
"00000111111110000111111110000000",
"00000011111111000111111110000000",
"00000011111111000111111110000000",
"00000011111111000111111100000000",
"00000011111111001111111100000000",
"00000011111111001111111100000000",
"00000011111111001111111100000000",
"00000001111111001111111100000000",
"00000001111111001111111100000000",
"00000001111111101111111000000000",
"00000001111111101111111000000000",
"00000001111111101111111000000000",
"00000001111111111111111000000000",
"00000000111111111111111000000000",
"00000000111111111111111000000000",
"00000000111111111111110000000000",
"00000000111111111111110000000000",
"00000000111111111111110000000000",
"00000000111111111111110000000000",
"00000000011111111111110000000000",
"00000000011111111111110000000000",
"00000000011111111111100000000000",
"00000000011111111111100000000000",
"00000000011111111111100000000000",
"00000000011111111111100000000000",
"00000000001111111111100000000000",
"00000000001111111111000000000000",
"00000000001111111111000000000000",
"00000000001111111111000000000000",
"00000000001111111111000000000000",
"00000000001111111111000000000000",
"00000000000111111111000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000010000111111111000",
"00111111111000010000111111111000",
"00111111111000111000111111111000",
"00111111111000111000111111111000",
"00111111111001111100111111111000",
"00111111111011111110111111111000",
"00111111111011111110111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111101111111111111000",
"00111111111111101111111111111000",
"00111111111111101111111111111000",
"00111111111111101111111111111000",
"00111111111111000111111111111000",
"00111111111111000111111111111000",
"00111111111111000111111111111000",
"00111111111111000111111111111000",
"00111111111110000011111111111000",
"00111111111110000011111111111000",
"00111111111110000011111111111000",
"00111111111110000011111111111000",
"00111111111100000001111111111000",
"00111111111100000001111111111000",
"00111111111100000001111111111000",
"00111111111100000001111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111111111111000000000000",
"00111111111111111111000000000000",
"00111111111111111111000000000000",
"00111111111111111111000000000000",
"00111111111111111111000000000000",
"00111111111111111111000000000000",
"00111111111111111111000000000000",
"00111111111111111111000000000000",
"00111111111111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111111111111111111100000",
"00011111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00011111111111111111111111110000",
"00011111111111111111111111110000",
"00000111111111111111111111000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111111111111111111100000",
"00011111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000011111111111111111000",
"00000000000011111111111111111000",
"00000000000011111111111111111000",
"00000000000011111111111111111000",
"00000000000011111111111111111000",
"00000000000011111111111111111000",
"00000000000011111111111111111000",
"00000000000011111111111111111000",
"00000000000011111111111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00011111111111111111111111110000",
"00011111111111111111111111110000",
"00000111111111111111111111000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111111111111111111100000",
"00011111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00011111111111111111111111110000",
"00011111111111111111111111110000",
"00000111111111111111111111000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111111111111111111111000",
"00011111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111111111111111111000000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111110000",
"00011111111111111111111111110000",
"00001111111111111111111111100000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111111111111111111000000",
"00011111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00011111111111111111111111110000",
"00011111111111111111111111100000",
"00000111111111111111111110000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111111111111111111100000",
"00011111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00011111111111111111111111111000",
"00001111111111111111111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111110000",
"00111111111111111111111111100000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000111111111111111111111000000",
"00001111111111111111111111100000",
"00011111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00011111111111111111111111110000",
"00001111111111111111111111100000",
"00000001111111111111111110000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000111111111111111111111111111",
"00001011111111111111111111111111",
"00001101111111111111111111111111",
"00001110111111111111111111111111",
"00001111000000000000000000000000",
"00001111001111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111100000000000001111",
"00001111011111100000000000000011",
"00001111011111100000000000000001",
"00001111011111100011111111100001",
"00001111011111100011111111110000",
"00001111011111100011111111111000",
"00001111011111100011111111111000",
"00001111011111100011111111111000",
"00001111011111100011111111110000",
"00001111011111100011111111100001",
"00001111011111100000000000000001",
"00001111011111100000000000000011",
"00001111011111100000000000001111",
"00001111011111100011111000011111",
"00001111011111100011111100001111",
"00001111011111100011111110000111",
"00001111011111100011111111000111",
"00001111011111100011111111000011",
"00001111011111100011111111100001",
"00001111011111100011111111110001",
"00001111011111100011111111110000",
"00001111011111100011111111111000",
"00001111011111100011111111111000",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111100111111111111111",
"00001111011111100111111111111111",
"00001111011111100111111111111111",
"00001111011111100111111100001100",
"00001111011111100111111000000100",
"00001111011111100111111001100100",
"00001111011111100111111000000100",
"00001111011111100111111001111110",
"00001111011111100111111001111110",
"00001111011111100000001000000111",
"00001111011111100000001100001111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111001111111111111111111111",
"00001111000000000000000000000000",
"00001110111111111111111111111111",
"00001101111111111111111111111111",
"00001011111111111111111111111111",
"00000111111111111111111111111111",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"11111111111111111111111111100000",
"11111111111111111111111111010000",
"11111111111111111111111110110000",
"11111111111111111111111101110000",
"00000000000000000000000011110000",
"11111111111111111111110011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111110011111111111011110000",
"11111111110011111111111011110000",
"11111111110011111111111011110000",
"11100001100000111111111011110000",
"11000000100000111111111011110000",
"11001100110011111111111011110000",
"11100111110011111111111011110000",
"11110001110011111111111011110000",
"11001000110011111111111011110000",
"11000000110000111111111011110000",
"01100001111000111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111110011111111011110000",
"11111111111110011111111011110000",
"11111111111110011111111011110000",
"11100110000110011111111011110000",
"11100100000010011111111011110000",
"11100100110010011111111011110000",
"01000100000010011111111011110000",
"01001100111110011111111011110000",
"00001100111110011111111011110000",
"00011100000010001111111011110000",
"10111110000110001111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111110011110000",
"00000000000000000000000011110000",
"11111111111111111111111101110000",
"11111111111111111111111110110000",
"11111111111111111111111111010000",
"11111111111111111111111111100000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000111111111111111111111111111",
"00001011111111111111111111111111",
"00001101111111111111111111111111",
"00001110111111111111111111111111",
"00001111000000000000000000000000",
"00001111001111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011110000000000000111111",
"00001111011110000000000000111111",
"00001111011110011111111111111111",
"00001111011110011111111111111111",
"00001111011110011111111111111100",
"00001111011110011111111111111000",
"00001111011110011111111111110001",
"00001111011110000000000001110011",
"00001111011110000000000001110001",
"00001111011110011111111111111000",
"00001111011110011111111111111100",
"00001111011110011111111111111111",
"00001111011110011111111111111111",
"00001111011110011111111111110011",
"00001111011110011111111111110001",
"00001111011110000000000000111000",
"00001111011110000000000000111100",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111100111110011111111",
"00001111011111100011100011111111",
"00001111011111100001000011111111",
"00001111011111100100010011000011",
"00001111011111100110110010000001",
"00001111011111100111110010011001",
"00001111011111100111110010000001",
"00001111011111100111110010011111",
"00001111011111100111110010011111",
"00001111011111100111110010000001",
"00001111011111100111110011000011",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111001111111111111111111111",
"00001111000000000000000000000000",
"00001110111111111111111111111111",
"00001101111111111111111111111111",
"00001011111111111111111111111111",
"00000111111111111111111111111111",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"11111111111111111111111111100000",
"11111111111111111111111111010000",
"11111111111111111111111110110000",
"11111111111111111111111101110000",
"00000000000000000000000011110000",
"11111111111111111111110011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"00001111111000001111111011110000",
"00000111110000000111111011110000",
"11100011100011100011111011110000",
"11110011000111110011111011110000",
"11111111001111111111111011110000",
"00011111001111111111111011110000",
"00000111001111111111111011110000",
"10000011001111111111111011110000",
"11110011001111111111111011110000",
"11110011000111110011111011110000",
"11100011100111100011111011110000",
"00000111110000000111111011110000",
"00001111111000001111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"00100011001110011111111011110000",
"00000001001110011111111011110000",
"00011001001110011111111011110000",
"00111001001110011111111011110000",
"00111001000110011111111011110000",
"00111001000000011111111011110000",
"00111001001000111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111110011110000",
"00000000000000000000000011110000",
"11111111111111111111111101110000",
"11111111111111111111111110110000",
"11111111111111111111111111010000",
"11111111111111111111111111100000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000010000000000000000",
"00000000000000011000000000000000",
"00000000000000011000000000000000",
"00000000000000111100000000000000",
"00000000000000111100000000000000",
"00000000000001111110000000000000",
"00000000000001111110000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000111111111100000000000",
"00000000000111111111100000000000",
"00000000001111111111110000000000",
"00000000001111111111110000000000",
"00000000011111111111111000000000",
"00000000011111111111111000000000",
"00000000111111111111111100000000",
"00000000111111111111111100000000",
"00000000111111111111111100000000",
"00000001111111111111111110000000",
"00000001111111111111111110000000",
"00000011111111111111111111000000",
"00000011111111111111111111000000",
"00000111111111111111111111100000",
"00000111111111111111111111100000",
"00001111111111111111111111110000",
"00001111111111111111111111110000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111111111111111111110000",
"00001111111111111111111111110000",
"00000111111111111111111111100000",
"00000111111111111111111111100000",
"00000011111111111111111111000000",
"00000011111111111111111111000000",
"00000001111111111111111110000000",
"00000001111111111111111110000000",
"00000000111111111111111100000000",
"00000000111111111111111100000000",
"00000000111111111111111100000000",
"00000000011111111111111000000000",
"00000000011111111111111000000000",
"00000000001111111111110000000000",
"00000000001111111111110000000000",
"00000000000111111111100000000000",
"00000000000111111111100000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000001111110000000000000",
"00000000000001111110000000000000",
"00000000000000111100000000000000",
"00000000000000111100000000000000",
"00000000000000011000000000000000",
"00000000000000011000000000000000",
"00000000000000010000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000111111111111111111111111111",
"00001011111111111111111111111111",
"00001101111111111111111111111111",
"00001110111111111111111111111111",
"00001111000000000000000000000000",
"00001111001111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111100000001111111111",
"00001111011111100000001111111111",
"00001111011111100111111111111110",
"00001111011111100111111111111110",
"00001111011111100000111001000111",
"00001111011111100000111000000011",
"00001111011111100111111000110011",
"00001111011111100111111001110011",
"00001111011111100111111001110011",
"00001111011111100000001001110011",
"00001111011111100000001001110011",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111101111111",
"00001111011111111111111001111111",
"00001111011111111111110001111111",
"00001111011111111111100001111111",
"00001111011111111111000000000000",
"00001111011111111110000000000000",
"00001111011111111111000000000000",
"00001111011111111111100001111111",
"00001111011111111111110001111111",
"00001111011111111111111001111111",
"00001111011111111111111101111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111011111111111111111111111",
"00001111001111111111111111111111",
"00001111000000000000000000000000",
"00001110111111111111111111111111",
"00001101111111111111111111111111",
"00001011111111111111111111111111",
"00000111111111111111111111111111",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"11111111111111111111111111100000",
"11111111111111111111111111010000",
"11111111111111111111111110110000",
"11111111111111111111111101110000",
"00000000000000000000000011110000",
"11111111111111111111110011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"00111111111111111111111011110000",
"00111111111111111111111011110000",
"00001111111111111111111011110000",
"00001100001100100111111011110000",
"00111000000100000111111011110000",
"00111001100100011111111011110000",
"00111000000100111111111011110000",
"00111001111100111111111011110000",
"00111001111100111111111011110000",
"00001000000100111111111011110000",
"10001100001100111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111000111111111111011110000",
"11111111000111111111111011110000",
"11111111000111111111111011110000",
"11111111000111111111111011110000",
"00000000000111111111111011110000",
"00000000000111111111111011110000",
"00000000000111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111111011110000",
"11111111111111111111110011110000",
"00000000000000000000000011110000",
"11111111111111111111111101110000",
"11111111111111111111111110110000",
"11111111111111111111111111010000",
"11111111111111111111111111100000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
others => (others => '1')
);

signal y_x : std_logic_vector(10 downto 0) := (others => '0');

begin

	y_x <= address_y & address_x;

	memory_read:process(clock)
	begin
		if(rising_edge(clock)) then
			if(read_enable = '1') then
				data_out <= rom(to_integer(unsigned(y_x)));
			end if;
		end if;
	end process;

end Behavioral;

