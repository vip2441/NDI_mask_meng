----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:40:14 10/22/2019 
-- Design Name: 
-- Module Name:    wall_obj - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity draw_arena is
    Port ( pix_x, pix_y : in  STD_LOGIC_VECTOR (10 downto 0);			--citace radku a sloupcu
           clk, enable : in  STD_LOGIC;						--hodiny pro rizeni procesu nacitani z pameti a signal pro aktivaci obvodu
			  obj_en: out std_logic;
           color : out  STD_LOGIC_vector(2 downto 0));		--vystupni barva
end draw_arena;


architecture Behavioral of draw_arena is

type ROM_type is array(0 to 4095) of std_logic_vector(2 downto 0);
constant rom : ROM_type := (

------------------------------------------zacatek steny--------------------------------------------------------
"001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "000", 
"111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", 
"111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", 
"111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", 
"111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "000", 
"111", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "000", 
"111", "111", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", 
"111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", 
"111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", 
"111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "001", "000", 
"111", "111", "111", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", 
"111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", 
"111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", 
"111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", 
"111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", 
"111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", 
"111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "001", "111", "001", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "111", "001", "111", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "111", "001", "111", "001", "111", "001", 
"111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", 
"111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", 
"111", "001", "111", "001", "111", "001", "111", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "111", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "111", "001", "111", "001", 
"111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", 
"111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", 
"111", "001", "111", "001", "111", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", 
"001", "111", "001", "111", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "111", "001", 
"111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", 
"111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", "111", "001", 
"111", "001", "111", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", 
"001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "000", "001", 
"000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", 
"000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", 
"000", "001", "000", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "000", "001", "000", 
"001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", 
"001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", 
"001", "000", "001", "000", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "000", "001", "000", "001", 
"000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", 
"000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", 
"000", "001", "000", "001", "000", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "000", "001", "000", "001", "000", 
"001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", 
"001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", 
"001", "000", "001", "000", "001", "000", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "001", "000", "001", "000", "001", "000", "001", 
"000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", 
"000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", 
"000", "001", "000", "001", "000", "001", "000", "001", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "001", "000", "001", "000", "001", "000", "001", "000", 
"001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", 
"001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", 
"001", "000", "001", "000", "001", "000", "001", "000", "001", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "111", "001", "000", "001", "000", "001", "000", "001", "000", "001", 
"000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", 
"000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", 
"000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "111", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", 
"001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", 
"001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", 
"001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "111", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", 
"000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", 
"000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", 
"000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "001", "001", "001", "000", 
"111", "111", "111", "111", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", 
"001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", 
"001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", 
"001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "001", "001", "000", 
"111", "111", "111", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", 
"000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", 
"000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", 
"000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "001", "000", 
"111", "111", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", 
"001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", 
"001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", 
"001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", 
"111", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", 
"000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", 
"000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", 
"000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "001", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000",
others => (others =>'0'));

signal cntx, cnty: natural range 0 to 1200 := 0;
constant dimm_x: natural range 0 to 800 := 512;				
constant dimm_y: natural range 0 to 600 := 448;

begin
	
	--pocitadla radku a sloupcu areny
	cntx <= to_integer(unsigned(pix_x));
	cnty <= to_integer(unsigned(pix_y));
	
	memory_driver: process(clk, enable, cntx, cnty)
	begin
		if(rising_edge(clk)) then
			if(enable = '1') then
				if(((cntx < 64 + dimm_x and cnty < 64) or
										(cntx < 64 and (cnty >= 64 and cnty < dimm_y)) or
										((cntx >=dimm_x and cntx < 64 + dimm_x) and (cnty >= 64 and cnty < dimm_y)) or
										(cntx < 64 + dimm_x and (cnty >= dimm_y and cnty < 64 + dimm_y)))) then
					obj_en <= '1';
					color <= rom(((cntx - dimm_x) mod 64)*64 + ((cnty - dimm_y) mod 64));
				elsif(cntx >= 64 and cntx < dimm_x and cnty >= 64 and cnty < dimm_y) then
					obj_en <= '1';
					color <= rom(((cntx - dimm_x) mod 64)*64 + ((cnty - dimm_y) mod 64) + 4096);
				else
					obj_en <= '0';
					color <= "000";
				end if;
			else
				obj_en <= '0';
				color <= "000";
			end if;
		end if;
	end process;
	
end Behavioral;

