----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:01:29 10/28/2019 
-- Design Name: 
-- Module Name:    graphic_rom - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity graphic_rom is
    Port ( clock, read_enable : in  STD_LOGIC;
           address_x: in  STD_LOGIC_VECTOR (11 downto 0);
			  address_y: in  STD_LOGIC_VECTOR (2 downto 0);
           data_out : out  STD_LOGIC_VECTOR (2 downto 0));
end graphic_rom;

architecture Behavioral of graphic_rom is

type ROM_type is array(0 to 32767) of std_logic_vector(2 downto 0);
constant rom : ROM_type := (
-----------------------------------------ZACATEK STENY-------------------------------------------------------
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", 
"111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "111", 
"111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "000", 
"000", "111", "000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", 
"111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "111", 
"111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "000", "000", "111", "000", 
"000", "111", "000", "000", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "000", "000", "111", "000", 
"000", "111", "000", "000", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "000", "000", "111", "000", 
"000", "111", "000", "000", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "000", "000", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "000", 
"000", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "000", "000", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "000", "000", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "000", 
"000", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "000", "000", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", 
"111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "111", 
"111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "000", 
"000", "111", "000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", 
"111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "111", 
"111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000",
---------------------------------------------KONEC STENY/ZACATEK PODLAHY-----------------------------------------
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "111", "000", "111", "000", 
"000", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "000", 
"000", "000", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "111", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "111", 
"000", "000", "000", "000", "000", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "000", "000", "000", "000", "111", "000", "000", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000",
-----------------------------------------------KONEC PODLAHY/ZACATEK KAMENU------------------------------------
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "111", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "000", "000", "000", "000", "111", "000", "111", "000", "111", "000", "000", "000", 
"000", "111", "111", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "000", "000", "000", "000", "111", "000", "111", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "111", "111", "000", "000", "000", 
"000", "111", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "111", "111", "111", "111", "000", "000", 
"000", "111", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "111", "111", "111", "111", "000", "000", 
"000", "111", "111", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "111", "111", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "000", "000", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "000", "000", "000", 
"000", "111", "000", "000", "000", "000", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", "000", 
"000", "111", "000", "000", "000", "000", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", "000", 
"000", "111", "111", "000", "000", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "111", "111", "000", "000", "000", 
"000", "111", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "111", "111", "111", "111", "000", "000", 
"000", "111", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "111", "111", "111", "111", "000", "000", 
"000", "111", "111", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "111", "111", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "000", "000", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "000", "000", "000", 
"000", "111", "000", "000", "000", "000", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", "000", 
"000", "111", "000", "000", "000", "000", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", "000", 
"000", "111", "111", "000", "000", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "000", "000", "000", "000", "111", "111", "111", "111", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "000", "000", "000", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000",
-----------------------------------------------KONEC KAMENU/ZACATEK HRACE-------------------------------------
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "111", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "111", "000", 
"000", "000", "000", "000", "000", "111", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "100", 
"100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", 
"110", "110", "110", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "000", "000", "100", 
"100", "100", "100", "100", "100", "100", "000", "000", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "000", "111", "000", "000", "110", "110", "110", "110", "110", 
"110", "110", "110", "000", "000", "100", "000", "100", "100", "100", "100", "100", "100", "000", "000", "000", 
"000", "100", "100", "100", "100", "100", "100", "100", "000", "000", "110", "110", "110", "110", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "100", "100", "100", 
"100", "111", "111", "111", "111", "100", "100", "100", "000", "000", "000", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "100", "100", "000", "100", "100", "100", "100", "100", "100", "000", "000", "000", 
"000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "000", "110", "110", "110", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "000", "111", "000", "100", "100", "100", "111", 
"111", "111", "111", "111", "111", "111", "100", "100", "100", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "000", "000", "100", "100", "000", "000", "100", "100", "100", "100", "100", "100", "000", "000", 
"000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "000", "110", "110", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "100", "100", "111", "111", 
"111", "111", "100", "100", "100", "100", "100", "100", "100", "000", "111", "000", "110", "110", "110", "110", 
"110", "110", "000", "000", "100", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "000", 
"000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "000", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "100", "100", "111", "111", "111", 
"111", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", 
"100", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "000", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "100", "111", "111", "111", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "100", "000", "000", "000", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "100", "100", "100", "100", "100", "000", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "000", "111", "000", "100", "111", "111", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "111", "000", "110", "110", 
"110", "110", "110", "000", "000", "000", "000", "000", "100", "100", "000", "000", "000", "000", "000", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "000", "000", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "110", "110", 
"110", "110", "110", "000", "000", "000", "000", "000", "100", "000", "000", "000", "000", "000", "100", "000", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "000", "000", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "100", "100", 
"000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "000", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "000", "000", "100", "100", "111", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "100", "100", "000", 
"000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "000", "000", "000", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "000", "000", "000", "100", "111", "111", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "111", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "100", "100", "000", 
"000", "000", "000", "000", "100", "100", "100", "000", "000", "000", "000", "000", "000", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "000", "111", "000", "100", "111", "111", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "100", "100", "100", "000", "000", "000", "100", "000", "000", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "000", "000", "100", "100", "111", "111", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "100", "100", "000", "000", "000", "000", "100", "000", "000", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "000", "000", "100", "100", "111", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "100", "000", "000", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "000", "000", "100", "100", "111", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "000", "111", "000", "110", "110", "110", "110", "110", 
"110", "110", "110", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "000", "000", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "000", "000", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "110", "110", "110", "110", "110", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "000", "000", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "000", "111", "000", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "000", "111", "000", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", "000", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "000", "000", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "100", "100", "100", "100", "000", 
"000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "111", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "111", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "111", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "111", "000", 
"111", "000", "111", "000", "000", "000", "000", "000", "000", "000", "111", "000", "111", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "110", "000", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "110", "000", "111", "000", "111", "000", "111", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "111", "000", 
"111", "000", "111", "000", "000", "000", "000", "000", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "111", "000", "111", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "111", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "111", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "100", "100", "100", "100", "000", 
"000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "000", "000", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "000", "111", "000", "100", "111", "111", "111", "111", "111", 
"111", "100", "100", "100", "000", "000", "000", "000", "000", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", "000", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "000", "000", "100", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "100", "100", "100", "000", "111", "000", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "000", "000", "100", "111", "111", "100", "100", "100", "100", 
"100", "100", "111", "111", "111", "100", "100", "000", "000", "000", "110", "110", "110", "110", "110", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "000", "000", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "111", "111", "111", "100", "100", "000", "000", "000", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "000", "000", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "111", "111", "111", "100", "000", "111", "000", "110", "110", "110", "110", "110", 
"110", "110", "110", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "000", "000", "100", "100", "111", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "111", "111", "111", "100", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "100", "000", "000", "110", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "000", "000", "100", "100", "111", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "100", "100", "000", "000", "000", "000", "100", "000", "000", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "000", "111", "000", "100", "111", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "100", "100", "100", "000", "000", "000", "100", "000", "000", "110", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "000", "000", "000", "100", "111", "111", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "111", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "100", "100", "000", 
"000", "000", "000", "000", "100", "100", "100", "000", "000", "000", "000", "000", "000", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "000", "000", "100", "111", "111", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "100", "100", "000", 
"000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "000", "000", "000", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "000", "000", "100", "100", "111", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "100", "100", 
"000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "000", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "000", "000", "100", "100", "111", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "110", "110", 
"110", "110", "110", "000", "000", "000", "000", "000", "100", "000", "000", "000", "000", "000", "100", "000", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "000", "111", "000", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "111", "000", "110", "110", 
"110", "110", "110", "000", "000", "000", "000", "000", "100", "100", "000", "000", "000", "000", "000", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "100", "000", "000", "000", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "100", "100", "100", "100", "100", "000", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", 
"100", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "000", "110", "110", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "111", "000", "110", "110", "110", "110", 
"110", "110", "000", "000", "100", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "000", 
"000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "000", "110", "110", "110", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "000", "111", "000", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "000", "000", "100", "100", "000", "000", "100", "100", "100", "100", "100", "100", "000", "000", 
"000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "000", "110", "110", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "100", "100", "000", "100", "100", "100", "100", "100", "100", "000", "000", "000", 
"000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "000", "110", "110", "110", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "000", "111", "000", "000", "110", "110", "110", "110", "110", 
"110", "110", "110", "000", "000", "100", "000", "100", "100", "100", "100", "100", "100", "000", "000", "000", 
"000", "100", "100", "100", "100", "100", "100", "100", "000", "000", "110", "110", "110", "110", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "100", 
"100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", 
"110", "110", "110", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "000", "000", "100", 
"100", "100", "100", "100", "100", "100", "000", "000", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "111", "000", 
"000", "000", "000", "000", "000", "111", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "111", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000",
---------------------------------------------KONEC HRACE/ZACATEK JIDLA-----------------------------------------
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "010", "010", "010", "010", 
"010", "010", "010", "010", "010", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "010", "110", "010", "110", "010", "010", "010", "010", "010", 
"010", "010", "010", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "010", "110", "010", "010", "010", 
"010", "010", "010", "010", "010", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "010", "110", "010", "110", "010", "010", "010", "010", 
"010", "010", "010", "010", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "010", "110", "010", "110", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "010", "110", "010", "110", "010", "010", "010", 
"010", "010", "010", "010", "010", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "010", "010", "110", "010", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "010", "010", "110", "010", "110", "010", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "010", "110", "010", "010", "010", "010", 
"010", "010", "010", "010", "010", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "010", "010", "110", "010", "110", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "010", "110", "010", "010", "010", 
"010", "010", "010", "010", "010", "010", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "010", "110", "010", "110", "010", "110", "010", 
"010", "010", "010", "010", "010", "010", "010", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "010", "110", "010", "010", 
"010", "010", "010", "010", "010", "010", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "010", "010", "110", "010", "110", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "010", "110", "010", "010", "010", 
"010", "010", "010", "010", "010", "010", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "010", "110", "010", "110", "010", "110", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "000", "000", "000", "110", "110", "110", "110", "110", "110", "010", "110", "010", "010", 
"010", "010", "010", "010", "010", "010", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "010", "010", "110", "010", "110", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "010", "010", "010", 
"010", "010", "010", "010", "010", "010", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "010", "010", "110", "010", "110", "010", "110", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "010", "110", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "010", "110", "010", "110", "010", "110", "010", "110", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "010", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "010", "010", "110", "010", "110", "010", "110", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "110", "000", "000", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "010", "110", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "010", "110", "010", "110", "010", "110", "010", "110", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "000", "000", "000", "000", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "010", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "010", "010", "110", "010", "110", "010", "110", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "000", "000", "000", "000", "000", "110", 
"110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "010", "110", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "010", "110", "010", "110", "010", "110", "010", "110", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "000", "000", "000", "110", "000", "000", "000", "000", "000", "110", "110", "010", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "010", "010", "110", "010", "110", "010", "110", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "010", "110", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "010", "110", "010", "110", "010", "110", "010", "110", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "010", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "010", "010", "110", "010", "110", "010", "110", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "010", "110", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "010", "110", "010", "110", "010", "110", "010", "110", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "010", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "010", "010", "110", "010", "110", "010", "110", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "000", "000", "000", "110", "000", "000", "000", "000", "000", "110", "010", "110", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "010", "110", "010", "110", "010", "110", "010", "110", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "000", "000", "000", "000", "000", "110", 
"110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "110", "010", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "010", "010", "110", "010", "110", "010", "110", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "000", "000", "000", "000", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "010", "110", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "010", "110", "010", "110", "010", "110", "010", "110", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "110", "000", "000", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "010", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "010", "010", "110", "010", "110", "010", "110", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "010", "110", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "010", "010", "110", "010", "110", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "010", "010", "010", 
"010", "010", "010", "010", "010", "010", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "010", "110", "010", "110", "010", "110", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "010", "110", "010", "010", 
"010", "010", "010", "010", "010", "010", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "010", "010", "110", "010", "110", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "000", "000", "000", "110", "110", "110", "110", "110", "010", "110", "010", "010", "010", 
"010", "010", "010", "010", "010", "010", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "010", "110", "010", "110", "010", "110", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "010", "110", "010", "010", 
"010", "010", "010", "010", "010", "010", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "010", "010", "110", "010", "110", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "010", "010", "010", "010", "010", "010", "010", "110", 
"110", "010", "110", "110", "110", "110", "110", "110", "110", "110", "110", "010", "110", "010", "010", "010", 
"010", "010", "010", "010", "010", "010", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "010", "010", "110", "010", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "010", "110", "010", "010", "010", "010", 
"010", "010", "010", "010", "010", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "010", "110", "010", "110", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "010", "110", "010", "110", "010", "010", "010", 
"010", "010", "010", "010", "010", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "010", "110", "010", "010", "010", 
"010", "010", "010", "010", "010", "010", "010", "010", "010", "010", "010", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "010", "110", "010", "110", "010", "010", "010", "010", 
"010", "010", "010", "010", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "010", "010", "010", "010", 
"010", "010", "010", "010", "010", "010", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "010", "110", "010", "110", "010", "010", "010", "010", "010", 
"010", "010", "010", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000",
others => (others => '0'));

signal y_x : std_logic_vector(14 downto 0) := (others => '0');

begin

	y_x <= address_y & address_x;

	memory_read:process(clock)
	begin
		if(falling_edge(clock)) then
			if(read_enable = '1') then
				data_out <= rom(to_integer(unsigned(y_x)));
			end if;
		end if;
	end process;

end Behavioral;

