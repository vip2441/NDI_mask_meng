----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:28:17 11/20/2019 
-- Design Name: 
-- Module Name:    gui_sprite_rom - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity gui_sprite_rom is
    Port ( clock, read_enable : in  STD_LOGIC;
           address_x: in  STD_LOGIC_VECTOR (10 downto 0);
			  address_y: in  STD_LOGIC_VECTOR (5 downto 0);
           data_out : out  STD_LOGIC_VECTOR (2 downto 0));
end gui_sprite_rom;

architecture Behavioral of gui_sprite_rom is

type ROM_type is array(0 to 131071) of std_logic_vector(2 downto 0);
constant rom : ROM_type := (
--Napis LEVEL
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000",
--Napis TAHY
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000",
--Tlacitko RESET
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", 
"111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", 
"111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "000", "000", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", "111", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", 
"111", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", "111", 
"111", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", "111", 
"111", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", 
"111", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", 
"111", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", "111", 
"111", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", "111", 
"111", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", "111", 
"111", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "111", "000", "000", "000", "000", 
"000", "000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", "111", 
"111", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "000", "000", "111", "111", "111", "111", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "111", 
"000", "000", "000", "000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "111", 
"111", "000", "000", "000", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "111", 
"111", "111", "000", "000", "000", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", "111", 
"111", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", "111", 
"111", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", 
"111", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", 
"111", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000",
--Tlacitko ENTER
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "000", "000", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "111", "111", "000", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "111", "111", "000", "111", "111", "000", "111", "111", "111", "111", "111", "111", "000", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "000", "000", "000", 
"000", "000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", 
"111", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "000", "000", "000", "000", 
"000", "000", "000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", 
"111", "111", "000", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", 
"111", "111", "000", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", 
"111", "111", "000", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", 
"000", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", 
"000", "000", "000", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"000", "000", "000", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "111", "111", "000", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"000", "000", "000", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "111", "111", "000", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", 
"000", "000", "000", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", 
"111", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", 
"111", "111", "000", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "000", "111", "111", "000", "111", "000", "111", "111", "111", "111", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "000", "000", "111", "111", "111", "000", "111", "111", "111", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", 
"000", "000", "000", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000",
--Tlacitko ESCAPE
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", 
"111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", 
"111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "000", "000", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "000", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "000", "000", "111", "111", "111", "111", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "000", "000", "111", "111", "111", "111", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "000", "000", "111", "111", "111", "111", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "111", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "000", "000", "111", "111", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "000", "000", "111", "111", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "000", "000", "111", "111", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "111", "000", "000", "000", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", "111", "111", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", "111", "111", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "000", "111", "111", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "111", "111", "111", "111", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "000", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "000", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000",
--Cislo NULA
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000",
--Cislo JEDNA
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000",
--Cislo DVA
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000",
--Cislo TRI
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000",
--Cislo CTYRI
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000",
--Cislo PET
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000",
--Cislo SEST
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000",
--Cislo SEDM
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000",
--Cislo OSM
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000",
--Cislo DEVET
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000",
--LOGO
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "100", "100", "000", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "100", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "100", "100", "000", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "100", "000", "000", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", 
"110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", 
"110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "100", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", "110", "110", "110", "110", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", "110", 
"110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", "110", 
"110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", "110", "110", "110", "110", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "100", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "110", "000", "110", "110", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", 
"110", "110", "110", "110", "110", "110", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", 
"100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "100", "100", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "100", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "100", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "100", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "100", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "100", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", 
"100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", 
"100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "100", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "100", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "100", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "100", "100", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "110", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "110", "110", "110", "110", 
"110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "110", "110", "110", "110", "110", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "110", "110", "110", "110", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", "110", "110", 
"110", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "110", "110", "110", "110", "110", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "110", "110", "110", "110", "110", "110", "000", "110", "000", "110", "000", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "110", 
"110", "110", "110", "110", "110", "000", "000", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "000", "110", "000", "110", "000", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "110", "110", "110", "110", "110", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "110", "000", "000", "000", "000", "000", "000", "000", "110", "000", "110", "000", "110", "000", "110", 
"110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "000", "110", "000", "110", "000", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "110", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", 
"000", "110", "000", "000", "000", "000", "000", "110", "110", "110", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", 
"111", "000", "000", "000", "000", "000", "000", "000", "110", "110", "000", "110", "000", "110", "000", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", 
"000", "110", "000", "000", "000", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", 
"111", "111", "000", "000", "000", "000", "000", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", 
"000", "110", "000", "000", "000", "110", "000", "110", "000", "000", "000", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", 
"111", "111", "111", "000", "000", "000", "000", "000", "110", "110", "000", "110", "000", "110", "000", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", 
"000", "110", "000", "000", "110", "000", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "111", "000", "000", "000", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "110", "000", "110", "000", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", 
"000", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", 
"000", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", 
"000", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "110", "000", "110", "000", "110", "000", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "110", "110", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", 
"000", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", 
"000", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "111", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", 
"000", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "110", "110", "000", "000", 
"000", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "110", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", 
"000", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "110", "110", "110", 
"111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "110", "110", "110", "110", "110", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"110", "110", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", 
"000", "110", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "110", "110", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", 
"110", "110", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "110", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "110", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", 
"100", "100", "110", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "110", "110", "000", "000", "000", "000", "110", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "110", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "110", "110", "110", "000", "000", "110", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "110", "110", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "000", "000", "000", "000", "110", "110", "110", "110", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "110", "000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "110", "110", "110", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "110", "000", "110", "000", "110", "000", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "100", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "000", 
"110", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "110", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "110", "110", "110", 
"000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "110", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "110", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "110", "110", "110", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "110", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "110", "110", "110", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "110", "110", "110", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "110", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "110", "000", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", 
"100", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "110", "000", "110", "000", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "000", "110", "000", "000", "000", "000", "000", "000", "000", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "110", "110", "000", "110", "000", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "110", "000", "110", "000", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "110", "110", "000", "110", "000", 
"110", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "110", "000", "110", "000", "110", 
"110", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", 
"000", "000", "000", "111", "110", "000", "000", "000", "000", "000", "110", "000", "110", "000", "000", "000", 
"000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "110", "110", "000", "110", "000", 
"110", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", 
"000", "000", "111", "111", "110", "000", "000", "000", "000", "110", "000", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "110", "000", "110", "000", "110", 
"110", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", 
"000", "111", "111", "111", "110", "000", "000", "000", "110", "000", "110", "000", "110", "000", "000", "000", 
"000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "110", "110", "000", "110", "000", 
"110", "000", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", 
"111", "111", "111", "000", "110", "000", "000", "110", "000", "110", "000", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "110", "000", "110", "000", "110", 
"110", "110", "110", "110", "110", "110", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "110", "000", "110", "000", "110", "000", "110", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "110", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "110", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "000", "000", "000", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "110", "000", "000", "000", "000", "000", "110", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "110", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "000", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "000", "000", "000", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "111", "111", "111", "111", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "110", "000", "000", "000", "000", "000", "110", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "111", "111", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", 
"000", "110", "000", "110", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "111", "110", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "110", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", 
"110", "000", "110", "000", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "111", "110", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "111", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "110", "000", "110", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"110", "000", "110", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"000", "110", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "111", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"110", "000", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "111", "111", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"000", "000", "000", "000", "000", "110", "000", "111", "111", "111", "111", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "000", "000", "000", "000", "110", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"111", "111", "111", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"000", "000", "000", "000", "000", "110", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "000", "000", "000", "000", "110", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "110", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"000", "000", "000", "000", "000", "110", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", "111", 
"111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "000", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", 
"111", "111", "111", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"000", "000", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", 
"000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "000", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", 
"000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", 
"110", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"000", "000", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", 
"000", "000", "000", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "000", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "110", "110", "110", "000", "110", "000", "110", "000", "110", "000", 
"000", "000", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "000", "000", "000", "000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "100", "100", "100", "110", "110", "110", "110", "000", "110", "000", "110", 
"000", "000", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "110", "110", "110", "110", "000", 
"000", "000", "000", "000", "000", "110", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "100", "000", "000", "000", 
"000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", "110", 
"000", "000", "000", "000", "000", "110", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "110", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "000", "000", "000", "000", "110", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"000", "000", "000", "000", "000", "110", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "110", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"110", "110", "110", "110", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "100", "100", "100", "100", "100", "100", "000", "100", "000", 
"000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "110", "110", "100", "100", "100", "100", "100", "100", "000", "100", 
"000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "110", "110", "100", "100", "100", "100", "100", "100", "000", 
"100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "000", "100", 
"000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "000", 
"100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "000", 
"100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"110", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"110", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"110", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", 
"100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"110", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", 
"100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"110", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "100", "100", "100", "100", "100", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "100", "100", "100", "100", "100", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "100", "100", "100", "100", "100", "110", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "100", "100", "100", "100", "100", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "100", "100", "100", "100", "100", "110", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "100", "100", "100", "100", "100", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "110", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "000", "000", "110", "000", "110", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "110", "110", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "110", "000", "110", "000", "110", "110", "110", "110", "110", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", 
"100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "110", "110", "110", "110", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", 
"100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "000", "110", "110", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "000", "000", "000", "000", "110", 
"110", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "110", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"000", "100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "000", 
"100", "000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"000", "100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "000", 
"100", "000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "000", "100", 
"000", "100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "000", 
"100", "000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "100", "100", "100", "100", "100", "000", "100", 
"000", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", 
"000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "000", "000", "000", "000", "000", "110", "110", "110", "000", "000", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "000", "000", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", 
"110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "111", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "110", "110", "110", "000", "000", "111", "111", "111", "000", "000", 
"110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", 
"110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "110", "110", "110", "110", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "100", "100", 
"100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "110", "110", "110", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "000", "000", "000", "000", "110", "110", "110", "110", "100", "100", "100", "100", "100", 
"100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "110", "110", "110", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "000", "000", "110", "110", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "110", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "100", "000", "000", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "100", "100", "000", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "000", "000", 
"000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "111", "100", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "111", "100", "100", "000", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "110", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "110", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", 
"110", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "000", "110", "000", "110", "000", "110", "000", "110", "000", "110", 
"000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "110", "000", "110", "000", "110", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "000", "110", "000", "110", "000", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "000", "000", "000", "000", "000", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "110", "000", "110", "000", "110", "000", "110", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", "000", "000", "000", "000", "000", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", "000", "000", "000", "000", "000", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "110", "000", "110", "000", "110", "000", "110", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", "000", "000", "000", "000", "000", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "110", "000", "110", "000", "110", "000", "110", "110", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", "000", "000", "000", "000", "000", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "110", "000", "110", "000", "110", "000", "110", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", "000", "000", "000", "000", "000", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "110", "000", "110", "000", "110", "000", "000", "110", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", "000", "000", "000", "000", "000", 
"000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "110", "000", "110", "000", "000", "000", "110", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", "000", "000", "000", "000", "000", 
"110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "110", "000", "110", "000", "000", "000", "000", "110", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "110", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "100", "110", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "100", "100", "100", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "000", "100", "000", "100", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "000", "100", "000", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "000", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "100", "100", "100", "100", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "000", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "100", "100", "100", "100", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "000", "000", "000", "000", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "100", "100", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"110", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "100", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"110", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "100", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"110", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "100", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"110", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"110", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", 
"100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"110", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", 
"100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"110", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"110", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "100", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "100", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "100", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "100", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "100", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "100", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "100", "100", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", 
"100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "100", "100", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", 
"100", "000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", "000", "100", 
"000", "100", "000", "100", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
others => (others => '0'));

signal y_x : std_logic_vector(16 downto 0) := (others => '0');

begin

	y_x <= address_y & address_x;

	memory_read:process(clock)
	begin
		if(rising_edge(clock)) then
			if(read_enable = '1') then
				data_out <= rom(to_integer(unsigned(y_x)));
			end if;
		end if;
	end process;
	
end Behavioral;

