----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:31:20 11/29/2019 
-- Design Name: 
-- Module Name:    ROM_lett_num - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ROM_lett_num is
	Port ( clock, read_enable : in  STD_LOGIC;
           address_x: in  STD_LOGIC_VECTOR (5 downto 0);
			  address_y: in  STD_LOGIC_VECTOR (4 downto 0);
           data_out : out  STD_LOGIC_VECTOR (0 to 31));
end ROM_lett_num;

architecture Behavioral of ROM_lett_num is

type ROM_type is array(0 to 2047) of std_logic_vector(0 to 31);
constant rom : ROM_type := (
	"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111111111111111111100000",
"00011111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111110000",
"00011111111111111111111111110000",
"00001111111111111111111111000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111111111111111111100000",
"00011111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111111111111111111000000",
"00111111111111111111111111000000",
"00111111111111111111111111000000",
"00111111111111111111111111000000",
"00111111111111111111111111000000",
"00111111111111111111111111000000",
"00111111111111111111111111000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111110000",
"00011111111111111111111111110000",
"00001111111111111111111111000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111000000000111111000000",
"00011111111000000000111111110000",
"00111111111100000000111111110000",
"00111111111100000000111111111000",
"00111111111100000000111111111000",
"00111111111110000000111111111000",
"00111111111110000000111111111000",
"00111111111110000000111111111000",
"00111111111111000000111111111000",
"00111111111111000000111111111000",
"00111111111111000000111111111000",
"00111111111111100000111111111000",
"00111111111111100000111111111000",
"00111111111111100000111111111000",
"00111111111111110000111111111000",
"00111111111111110000111111111000",
"00111111111111110000111111111000",
"00111111111111111000111111111000",
"00111111111111111000111111111000",
"00111111111111111000111111111000",
"00111111111111111100111111111000",
"00111111111111111100111111111000",
"00111111111111111100111111111000",
"00111111111111111110111111111000",
"00111111111111111110111111111000",
"00111111111111111110111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111011111111111111111000",
"00111111111011111111111111111000",
"00111111111011111111111111111000",
"00111111111001111111111111111000",
"00111111111001111111111111111000",
"00111111111000111111111111111000",
"00111111111000111111111111111000",
"00111111111000111111111111111000",
"00111111111000011111111111111000",
"00111111111000011111111111111000",
"00111111111000011111111111111000",
"00111111111000001111111111111000",
"00111111111000001111111111111000",
"00111111111000000111111111111000",
"00111111111000000111111111111000",
"00111111111000000111111111111000",
"00111111111000000011111111111000",
"00111111111000000011111111111000",
"00111111111000000011111111111000",
"00111111111000000001111111111000",
"00111111111000000001111111111000",
"00111111111000000000111111111000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111111111111111111100000",
"00111111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111110000",
"00111111111111111111111111100000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111111111111111111000000",
"00111111111111111111111111100000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111100000",
"00111111111111111111111111000000",
"00111111111000111111110000000000",
"00111111111000111111110000000000",
"00111111111000111111111000000000",
"00111111111000011111111000000000",
"00111111111000011111111000000000",
"00111111111000011111111100000000",
"00111111111000001111111100000000",
"00111111111000001111111110000000",
"00111111111000000111111110000000",
"00111111111000000111111110000000",
"00111111111000000111111111000000",
"00111111111000000011111111000000",
"00111111111000000011111111100000",
"00111111111000000011111111100000",
"00111111111000000001111111110000",
"00111111111000000001111111110000",
"00111111111000000000111111110000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000011111111100",
"00111111111000000000011111111100",
"00111111111000000000011111111110",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111110000000111111111000",
"00011111111111000000111111111000",
"00011111111111000000111111111000",
"00001111111111000000111111111000",
"00001111111111100000111111111000",
"00000111111111100000111111111000",
"00000111111111110000111111111000",
"00000011111111110000111111111000",
"00000011111111111000111111111000",
"00000011111111111000000000000000",
"00000001111111111100000000000000",
"00000001111111111100000000000000",
"00000000111111111110000000000000",
"00000000111111111110000000000000",
"00000000011111111111000000000000",
"00000000011111111111000000000000",
"00000000001111111111000000000000",
"00000000001111111111100000000000",
"00000000000111111111100000000000",
"00000000000111111111110000000000",
"00000000000011111111110000000000",
"00000000000011111111111000000000",
"00000000000001111111111000000000",
"00000000000001111111111100000000",
"00000000000000111111111100000000",
"00000000000000111111111110000000",
"00111111111000011111111110000000",
"00111111111000011111111110000000",
"00111111111000011111111111000000",
"00111111111000001111111111000000",
"00111111111000001111111111100000",
"00111111111000000111111111100000",
"00111111111000000111111111110000",
"00111111111000000011111111110000",
"00111111111000000011111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111111111111111111111110",
"00111111111111111111111111111110",
"00111111111111111111111111111110",
"00111111111111111111111111111110",
"00111111111111111111111111111110",
"00111111111111111111111111111110",
"00111111111111111111111111111110",
"00111111111111111111111111111110",
"00111111111111111111111111111110",
"00111111111000011111111100000000",
"00111111111000011111111100000000",
"00111111111000011111111100000000",
"00111111111000011111111100000000",
"00111111111000011111111100000000",
"00111111111000011111111100000000",
"00111111111000011111111100000000",
"00111111111000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000011111111100000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111000000000111111110000",
"00111111111000000001111111110000",
"00111111111000000001111111110000",
"00111111111000000001111111110000",
"00011111111000000001111111110000",
"00011111111000000001111111110000",
"00011111111100000001111111100000",
"00011111111100000001111111100000",
"00011111111100000001111111100000",
"00011111111100000011111111100000",
"00001111111100000011111111100000",
"00001111111100000011111111100000",
"00001111111100000011111111000000",
"00001111111100000011111111000000",
"00001111111110000011111111000000",
"00001111111110000011111111000000",
"00000111111110000011111111000000",
"00000111111110000111111111000000",
"00000111111110000111111110000000",
"00000111111110000111111110000000",
"00000111111110000111111110000000",
"00000111111110000111111110000000",
"00000011111111000111111110000000",
"00000011111111000111111110000000",
"00000011111111000111111100000000",
"00000011111111001111111100000000",
"00000011111111001111111100000000",
"00000011111111001111111100000000",
"00000001111111001111111100000000",
"00000001111111001111111100000000",
"00000001111111101111111000000000",
"00000001111111101111111000000000",
"00000001111111101111111000000000",
"00000001111111111111111000000000",
"00000000111111111111111000000000",
"00000000111111111111111000000000",
"00000000111111111111110000000000",
"00000000111111111111110000000000",
"00000000111111111111110000000000",
"00000000111111111111110000000000",
"00000000011111111111110000000000",
"00000000011111111111110000000000",
"00000000011111111111100000000000",
"00000000011111111111100000000000",
"00000000011111111111100000000000",
"00000000011111111111100000000000",
"00000000001111111111100000000000",
"00000000001111111111000000000000",
"00000000001111111111000000000000",
"00000000001111111111000000000000",
"00000000001111111111000000000000",
"00000000001111111111000000000000",
"00000000000111111111000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000010000111111111000",
"00111111111000010000111111111000",
"00111111111000111000111111111000",
"00111111111000111000111111111000",
"00111111111001111100111111111000",
"00111111111011111110111111111000",
"00111111111011111110111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111101111111111111000",
"00111111111111101111111111111000",
"00111111111111101111111111111000",
"00111111111111101111111111111000",
"00111111111111000111111111111000",
"00111111111111000111111111111000",
"00111111111111000111111111111000",
"00111111111111000111111111111000",
"00111111111110000011111111111000",
"00111111111110000011111111111000",
"00111111111110000011111111111000",
"00111111111110000011111111111000",
"00111111111100000001111111111000",
"00111111111100000001111111111000",
"00111111111100000001111111111000",
"00111111111100000001111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000111111100000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111111111111000000000000",
"00111111111111111111000000000000",
"00111111111111111111000000000000",
"00111111111111111111000000000000",
"00111111111111111111000000000000",
"00111111111111111111000000000000",
"00111111111111111111000000000000",
"00111111111111111111000000000000",
"00111111111111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00000000000111111111000000000000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111111111111111111100000",
"00011111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00011111111111111111111111110000",
"00011111111111111111111111110000",
"00000111111111111111111111000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111111111111111111100000",
"00011111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000011111111111111111000",
"00000000000011111111111111111000",
"00000000000011111111111111111000",
"00000000000011111111111111111000",
"00000000000011111111111111111000",
"00000000000011111111111111111000",
"00000000000011111111111111111000",
"00000000000011111111111111111000",
"00000000000011111111111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00011111111111111111111111110000",
"00011111111111111111111111110000",
"00000111111111111111111111000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111111111111111111100000",
"00011111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00011111111111111111111111110000",
"00011111111111111111111111110000",
"00000111111111111111111111000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111111111111111111111000",
"00011111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111000000000000000000000",
"00111111111111111111111111000000",
"00111111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111110000",
"00011111111111111111111111110000",
"00001111111111111111111111100000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111111111111111111000000",
"00011111111111111111111111110000",
"00111111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00011111111111111111111111110000",
"00011111111111111111111111100000",
"00000111111111111111111110000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111111111111111111100000",
"00011111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00011111111111111111111111111000",
"00001111111111111111111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00000000000000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111110000",
"00111111111111111111111111100000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000111111111111111111111000000",
"00001111111111111111111111100000",
"00011111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111000000000111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00111111111111111111111111111000",
"00011111111111111111111111110000",
"00001111111111111111111111100000",
"00000001111111111111111110000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"10111111111111111111111111111111",
"11111111111111111111111111111110",
"01011111111111111111111111111111",
"11111111111111111111111111111100",
"10101111111111111111111111111111",
"11111111111111111111111111111000",
"01010111111111111111111111111111",
"11111111111111111111111111110000",
"10101011111111111111111111111111",
"11111111111111111111111111100000",
"01010101111111111111111111111111",
"11111111111111111111111111000000",
"10101010111111111111111111111111",
"11111111111111111111111110000000",
"01010101011000000000000000000000",
"00000000000000000000000000000000",
"10101010100111111111111111111111",
"11111111111111111111100000000000",
"01010101001111111111111111111111",
"11111111111111111111110000000000",
"10101010011111111111111111111111",
"11111111111111111111111000000000",
"01010100111111111111111111111111",
"11111111111111111111111100000000",
"10101010111111111111111111111111",
"11111111111111111111111100000000",
"01010100111111111111111111111111",
"11111111111111111111111100000000",
"10101010111111111111111111111111",
"11111111111111111111111100000000",
"01010100111111111111111100000000",
"00001111111111111111111100000000",
"10101010111111111111111100000000",
"00000011111111111111111100000000",
"01010100111111111111111100000000",
"00000001111111111111111100000000",
"10101010111111111111111100001111",
"11000001111111111111111100000000",
"01010100111111111111111100001111",
"11100001111111111111111100000000",
"10101010111111111111111100001111",
"11100001111111111111111100000000",
"01010100111111111111111100001111",
"11100001111111111111111100000000",
"10101010111111111111111100001111",
"11100001111111111111111100000000",
"01010100111111111111111100001111",
"11000001111111111111111100000000",
"10101010111111111111111100000000",
"00000001111111111111111100000000",
"01010100111111111111111100000000",
"00000001111111111111111100000000",
"10101010111111111111111100000000",
"00000011111111111111111100000000",
"01010100111111111111111100000000",
"01111111111111111111111100000000",
"10101010111111111111111100001000",
"00111111111111111111111100000000",
"01010100111111111111111100001000",
"00111111111111111111111100000000",
"10101010111111111111111100001100",
"00011111111111111111111100000000",
"01010100111111111111111100001110",
"00011111111111111111111100000000",
"10101010111111111111111100001111",
"00001111111111111111111100000000",
"01010100111111111111111100001111",
"00000111111111111111111100000000",
"10101010111111111111111100001111",
"10000011111111111111111100000000",
"01010100111111111111111100001111",
"11000001111111111111111100000000",
"10101010111111111111111100001111",
"11000001111111111111111100000000",
"01010100111111111111111111111111",
"11111111111111111111111100000000",
"10101010111111111111111111111111",
"11111111111111111111111100000000",
"01010100111111111111111111111111",
"11111111111111111111111100000000",
"10101010111111111111111111111111",
"11111111111111111111111100000000",
"01010100111111111111111111111111",
"11111111111111111111111100000000",
"10101010111111111111111111111111",
"11111111111111111111111100000000",
"01010100111111111000011000001100",
"00110000010000011111111100000000",
"10101010111111111011101011111011",
"11010111111101111111111100000000",
"01010100111111111011101011111011",
"11110111111101111111111100000000",
"10101010111111111000011000111100",
"00110001111101111111111100000000",
"01010100111111111010111011111111",
"11010111111101111111111100000000",
"10101010111111111011011011111011",
"11010111111101111111111100000000",
"01010100111111111011101000001100",
"00110000011101111111111100000000",
"10101010111111111111111111111111",
"11111111111111111111111100000000",
"01010100111111111111111111111111",
"11111111111111111111111100000000",
"10101010111111111111111111111111",
"11111111111111111111111100000000",
"01010100011111111111111111111111",
"11111111111111111111111000000000",
"10101010001111111111111111111111",
"11111111111111111111110000000000",
"01010100000111111111111111111111",
"11111111111111111111100000000000",
"10101010000000000000000000000000",
"00000000000000000000000000000000",
"01010100000000000000000000000000",
"00000000000000000000000000000000",
"10101000000000000000000000000000",
"00000000000000000000000000000000",
"01010000000000000000000000000000",
"00000000000000000000000000000000",
"10100000000000000000000000000000",
"00000000000000000000000000000000",
"01000000000000000000000000000000",
"00000000000000000000000000000000",
"10000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"10111111111111111111111111111111",
"11111111111111111111111111111110",
"01011111111111111111111111111111",
"11111111111111111111111111111100",
"10101111111111111111111111111111",
"11111111111111111111111111111000",
"01010111111111111111111111111111",
"11111111111111111111111111110000",
"10101011111111111111111111111111",
"11111111111111111111111111100000",
"01010101111111111111111111111111",
"11111111111111111111111111000000",
"10101010111111111111111111111111",
"11111111111111111111111110000000",
"01010101011000000000000000000000",
"00000000000000000000000000000000",
"10101010100111111111111111111111",
"11111111111111111111100000000000",
"01010101001111111111111111111111",
"11111111111111111111110000000000",
"10101010011111111111111111111111",
"11111111111111111111111000000000",
"01010100111111111111111111111111",
"11111111111111111111111100000000",
"10101010111111111111111111111111",
"11111111111111111111111100000000",
"01010100111111111111111111111111",
"11111111111111111111111100000000",
"10101010111111111111111111111111",
"11111111111111111111111100000000",
"01010100111111111111111111111111",
"11111111111111111111111100000000",
"10101010111111111111111111111111",
"11111111111111111111111100000000",
"01010100111111111111111111111111",
"11111111111111111111111100000000",
"10101010111111111111111111111111",
"11111111111111111111111100000000",
"01010100111111111111111111111111",
"11111111111111111111111100000000",
"10101010111111111111111111111111",
"11111111111111111111111100000000",
"01010100111111111111000000001111",
"11111111111111111111111100000000",
"10101010111111111111000000001111",
"11111111111111111111111100000000",
"01010100111111111111001111111111",
"11111111111111111111111100000000",
"10101010111111111111001111111100",
"00011100000111111111111100000000",
"01010100111111111111001111111000",
"00001000000011111111111100000000",
"10101010111111111111000001111001",
"11001001110011111111111100000000",
"01010100111111111111000001111001",
"11111001111111111111111100000000",
"10101010111111111111001111111000",
"00011001111111111111111100000000",
"01010100111111111111001111111100",
"00001001111111111111111100000000",
"10101010111111111111001111111111",
"11001001111111111111111100000000",
"01010100111111111111001111111001",
"11001001110011111111111100000000",
"10101010111111111111000000001000",
"00001000000011111111111100000000",
"01010100111111111111000000001100",
"00011100000111111111111100000000",
"10101010111111111111111111111111",
"11111111111111111111111100000000",
"01010100111111111111111111111111",
"11111111111111111111111100000000",
"10101010111111111111111111111111",
"11111111111111111111111100000000",
"01010100111111111111111111111111",
"11111111111111111111111100000000",
"10101010111111111111111111111111",
"11111111111111111111111100000000",
"01010100111111111111111111111111",
"11111111111111111111111100000000",
"10101010111111111111111111111111",
"11111111111111111111111100000000",
"01010100111111111111111111111111",
"11111111111111111111111100000000",
"10101010111111111101110110001101",
"11010000011000111111111100000000",
"01010100111111111101101101110100",
"11010111110111011111111100000000",
"10101010111111111101011101110101",
"01010111110111111111111100000000",
"01010100111111111100111101110101",
"01010000110111111111111100000000",
"10101010111111111101011101110101",
"10010111110111111111111100000000",
"01010100111111111101101101110101",
"11010111110111011111111100000000",
"10101010111111111101110110001101",
"11010000011000111111111100000000",
"01010100111111111111111111111111",
"11111111111111111111111100000000",
"10101010111111111111111111111111",
"11111111111111111111111100000000",
"01010100111111111111111111111111",
"11111111111111111111111100000000",
"10101010111111111111111111111111",
"11111111111111111111111100000000",
"01010100011111111111111111111111",
"11111111111111111111111000000000",
"10101010001111111111111111111111",
"11111111111111111111110000000000",
"01010100000111111111111111111111",
"11111111111111111111100000000000",
"10101010000000000000000000000000",
"00000000000000000000000000000000",
"01010100000000000000000000000000",
"00000000000000000000000000000000",
"10101000000000000000000000000000",
"00000000000000000000000000000000",
"01010000000000000000000000000000",
"00000000000000000000000000000000",
"10100000000000000000000000000000",
"00000000000000000000000000000000",
"01000000000000000000000000000000",
"00000000000000000000000000000000",
"10000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",

others => (others => '1')
);

signal y_x : std_logic_vector(10 downto 0) := (others => '0');

begin

	y_x <= address_y & address_x;

	memory_read:process(clock)
	begin
		if(rising_edge(clock)) then
			if(read_enable = '1') then
				data_out <= rom(to_integer(unsigned(y_x)));
			end if;
		end if;
	end process;

end Behavioral;

