----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:03:29 11/04/2019 
-- Design Name: 
-- Module Name:    stone_obj - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity stone_obj is
    Port ( pix_x, pix_y : in  STD_LOGIC_VECTOR (10 downto 0);
           enable, clk : in  STD_LOGIC;
           color : out  STD_LOGIC_VECTOR (2 downto 0));
end stone_obj;

architecture Behavioral of stone_obj is

type ROM_type is array(0 to 4095) of std_logic_vector(2 downto 0);
constant rom : ROM_type := (
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", 
"000", "111", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "000", "000", "000", "000", "111", "000", "111", "000", "111", "000", "000", "000", 
"000", "111", "111", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "000", "000", "000", "000", "111", "000", "111", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "000", "000", "111", "000", "111", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", 
"000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "111", "000", 
"111", "000", "111", "000", "111", "000", "111", "000", "111", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "111", "111", "000", "000", "000", 
"000", "111", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "111", "111", "111", "111", "000", "000", 
"000", "111", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "111", "111", "111", "111", "000", "000", 
"000", "111", "111", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "111", "111", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "000", "000", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "000", "000", "000", 
"000", "111", "000", "000", "000", "000", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", "000", 
"000", "111", "000", "000", "000", "000", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", "000", 
"000", "111", "111", "000", "000", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "111", "111", "000", "000", "000", 
"000", "111", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "111", "111", "111", "111", "000", "000", 
"000", "111", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "111", "111", "111", "111", "000", "000", 
"000", "111", "111", "000", "000", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "111", "111", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "000", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "000", "000", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "000", "000", "000", 
"000", "111", "000", "000", "000", "000", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", "000", 
"000", "111", "000", "000", "000", "000", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", "000", 
"000", "111", "111", "000", "000", "111", "111", "111", "110", "110", "110", "110", "110", "110", "110", "110", 
"110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "111", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "111", "000", "000", "000", "000", "111", "111", "111", "111", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "111", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "111", "111", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "111", "000", "000", "000", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", 
"000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000");

signal cntx, cnty: integer := 0;

begin

	cntx <= to_integer(unsigned(pix_x));
	cnty <= to_integer(unsigned(pix_y));
	
	process(clk,cntx, cnty, enable)
	begin
		if(rising_edge(clk)) then
			if(enable = '1') then
				color <= rom((cntx mod 64)*64 + (cnty mod 64));
			else
				color <= "000";
			end if;
		end if;
	end process;


end Behavioral;

