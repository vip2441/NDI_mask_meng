----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:16:17 11/28/2019 
-- Design Name: 
-- Module Name:    sprite_grayscale_ROM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity sprite_grayscale_ROM is
	Port ( clock, read_enable : in  STD_LOGIC;
           addr: in  STD_LOGIC_VECTOR (7 downto 0);
           data_out : out  STD_LOGIC_VECTOR (0 to 31));
end sprite_grayscale_ROM;

architecture Behavioral of sprite_grayscale_ROM is

	type ROM_type is array(0 to 255) of std_logic_vector(0 to 31);
	constant rom : ROM_type := (
	"00000000000000000000000000000000","00000000000000000000000000000000",
	"01111111111111111111111111111111","11111111111111111111111111111110",
	"01001111111100111111110011111111","00111111100111111110011111110010",
	"01001111111100111111110011111111","00111111100111111110011111110010",
	"01111111111111111111111111111111","11111111111111111111111111111110",
	"01111000000000000000000000000000","00000000000000000000000000011110",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01001010101010101010101010101010","10101010101010101010101010010010",
	"01001001010101010101010101010101","01010101010101010101010101010010",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01001010101010101010101010101010","10101010101010101010101010010010",
	"01001001010101010101010101010101","01010101010101010101010101010010",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01001010101010101010101010101010","10101010101010101010101010010010",
	"01001001010101010101010101010101","01010101010101010101010101010010",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01001001010101010101010101010101","01010101010101010101010101010010",
	"01001010101010101010101010101010","10101010101010101010101010010010",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01001001010101010101010101010101","01010101010101010101010101010010",
	"01001010101010101010101010101010","10101010101010101010101010010010",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01111010101010101010101010101010","10101010101010101010101010011110",
	"01111001010101010101010101010101","01010101010101010101010101011110",
	"01111000000000000000000000000000","00000000000000000000000000011110",
	"01111111111111111111111111111111","11111111111111111111111111111110",
	"01001111111100111111110011111111","00111111100111111110011111110010",
	"01001111111100111111110011111111","00111111100111111110011111110010",
	"01111111111111111111111111111111","11111111111111111111111111111110",
	"00000000000000000000000000000000","00000000000000000000000000000000",
	------------------------------konec steny/zacatek podlahy------------
	"00000000000000000000000000000000","00000000000000000000000000000000",
	"01010101010101010101010101010101","01010101010101010101010101010100",
	"00101010101010101010101010101010","10101010101010101010101010101010",
	"01010101010101010101010101010101","01010101010101010101010101010100",
	"00101010101010101010101010101010","10101010101010101010101010100000",
	"01010101010101010101010101010101","01010101010101010101010101000100",
	"00101010101010101010101010101010","10101010101010101010101010001010",
	"01010101010101010101010101010101","01010101010101010101010101000100",
	"00101010101010101010101010101010","10101010101010101010101010001010",
	"01010101010101010101010101010101","01010101010101010101010100010100",
	"00101010101010101010101010101010","10101010101000000010101000001010",
	"00010101010101010101010101010101","01010101010000000000010100010100",
	"00001010101010101010101010101010","10101010100000100000000000101010",
	"01000101010101010001010101010101","01010101000101010000000101010100",
	"00100010101010000010101010101010","10101010101010101010001010101010",
	"01010001010100000101010101010101","01010101010101010100010101010100",
	"00101000001000101010101010101010","10101010101010101010001010101010",
	"01010100000000010101010101010101","01010101010101010100010101010100",
	"00101010000000101010101010101010","10101010101010101000101010101010",
	"01010101010000010101010101010101","01010101010101000001010101010100",
	"00101010101010001010101010101010","10101010101010100010101010101010",
	"01010101010101000101010101010101","01010101010101000101010101010100",
	"00101010101010101010101010101010","10101010101010001010101010101010",
	"01010101010101000101010101010101","01010101010101010101010101010100",
	"00101010101010101010101010101010","10101010101010101010101010101010",
	"01010101010101010101010101010101","01010101010101010101010101010100",
	"00101010101010101010101010101010","10101010101010101010101010101010",
	"01010101010101010101010101010101","01010101010101010101010101010100",
	"00101010101010101010101010101010","10101010101010101010101010101010",
	"01010101010101010101010101010101","01010101010101010101010101010100",
	"00101010101010101010101010101010","10101010101010101010101010101010",
	"01010101010101010101010101010101","01010101010101010101010101010100",
	"00101010101010101010101010101010","10101010101010101010101010101010",
	"01010101010101010101010101010101","01010101010101010101010101010100",
	"00101010101010101010101010101010","10101010101010101010101010101010",
	"01010101010101010101010101010101","01010101010101010101010101010100",
	"00101010101010101010101010101010","10101010101010101010101010101010",
	"01010101010101010101010101010101","01010101010101010101010101010100",
	"00101010101010101010101010101010","10101010101010101010101010101010",
	"01010101010101010101010101010101","01010101010101010101010101010100",
	"00101010101010101010101010101010","10101010101010101010101010101010",
	"01010101010101010101010101010101","01010101010101010101010101010100",
	"00101010101010101010101010101010","10101010101010101010101010101010",
	"01010101010101010101010101010101","01010101010101010101010101010100",
	"00101010101010101010101010101010","10101010101010101010101010101010",
	"01010101010101010101010101010101","01010101010101010101010101010100",
	"00101010101010101010101010101010","10101010101010101010101010101010",
	"01010101010101010101010101010101","01010101010101010101010101010100",
	"00101010101010101010101010101010","10101010101010101010101010101010",
	"01010101010101010101010101010101","01010101010101010101010101010100",
	"00101010101010101010101010101010","10101010101010101010101010100000",
	"01010101010101010101010101010101","01010101010101010101010101000000",
	"00101010101010101010101010101010","10101010101010101010101010001010",
	"01010101010101010101010101010101","01010101010101010101010100010100",
	"00000010101010101010101010101000","10101010101010101000000000101010",
	"01010001010101010101010101010001","01010101010101010101000101010100",
	"00101010101010101010101010100010","10101010101010101010101010101010",
	"01010101010101010101010101000101","01010101010101010101010101010100",
	"00101010101010101010101010001010","10101010101010101010101010101010",
	"01010101010101010101010101000101","01010101010101010101010101010100",
	"00101010101010101010101010001010","10101010101010101010101010101010",
	"01010101010101010101010101010101","01010101010101010101010101010100",
	"00101010101010101010101010001010","10101010101010101010101010101010",
	"00000000000000000000000000000000","00000000000000000000000000000000"
	--------------------------konec podlahy/zacatek neceho----------------
	);

begin
	
	memory_read:process(clock)
	begin
		if(rising_edge(clock)) then
			if(read_enable = '1') then
				data_out <= rom(to_integer(unsigned(addr)));
			end if;
		end if;
	end process;


end Behavioral;

