----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:01:29 10/28/2019 
-- Design Name: 
-- Module Name:    graphic_rom - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity graphic_rom is
    Port ( clock, we, en: in  STD_LOGIC;
				data_in: in std_logic_vector(1 downto 0);
           address_x1, address_x2: in  STD_LOGIC_VECTOR (11 downto 0);
			  address_y1, address_y2: in  STD_LOGIC_VECTOR (3 downto 0);
           data_out1, data_out2 : out  STD_LOGIC_VECTOR (1 downto 0));
end graphic_rom;

architecture Behavioral of graphic_rom is

type ROM_type is array(0 to 65535) of std_logic_vector(1 downto 0);
signal rom : ROM_type := (
-------------------------------------------ZACATEK STENY--------------------------------------------------------------
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00",
"00","01","00","00","01","01","01","01","01","01","01","01","00","00","01","01","01","01","01","01","01","01","00","00","01","01","01","01","01","01","01","01",
"00","00","01","01","01","01","01","01","01","00","00","01","01","01","01","01","01","01","01","00","00","01","01","01","01","01","01","01","00","00","01","00",
"00","01","00","00","01","01","01","01","01","01","01","01","00","00","01","01","01","01","01","01","01","01","00","00","01","01","01","01","01","01","01","01",
"00","00","01","01","01","01","01","01","01","00","00","01","01","01","01","01","01","01","01","00","00","01","01","01","01","01","01","01","00","00","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00",
"00","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","01","01","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","00","00","01","00",
"00","01","00","00","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","00","00","01","00",
"00","01","00","00","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","00","00","01","00",
"00","01","00","00","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","00","00","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","00",
"00","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","00","00","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","00","00","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","00",
"00","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","00","00","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","01","01","01","01","00",
"00","01","01","01","01","00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","01","01","01","00",
"00","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00",
"00","01","00","00","01","01","01","01","01","01","01","01","00","00","01","01","01","01","01","01","01","01","00","00","01","01","01","01","01","01","01","01",
"00","00","01","01","01","01","01","01","01","00","00","01","01","01","01","01","01","01","01","00","00","01","01","01","01","01","01","01","00","00","01","00",
"00","01","00","00","01","01","01","01","01","01","01","01","00","00","01","01","01","01","01","01","01","01","00","00","01","01","01","01","01","01","01","01",
"00","00","01","01","01","01","01","01","01","00","00","01","01","01","01","01","01","01","01","00","00","01","01","01","01","01","01","01","00","00","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
--------------------------------------------KONEC STENY/ZACATEK PODLAHY-----------------------------------------------------------
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
-------------------------------------------KONEC PODLAHY/ZACATEK KAMENU----------------------------------------------------
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"00","01","00","01","00","01","00","01","00","00","00","01","00","01","00","01","00","01","00","01","00","01","00","00","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","00","00","01","00","01","00","01","00","01","00","01","00","01","00","00","00","01","00","01","00","01","00","01","00","00",
"00","01","01","00","01","00","01","00","00","00","00","00","01","00","01","00","01","00","01","00","01","00","00","00","00","00","01","00","01","00","01","00",
"01","00","01","00","01","00","00","00","00","00","01","00","01","00","01","00","01","00","01","00","00","00","00","00","01","00","01","00","01","00","00","00",
"00","01","01","01","00","01","00","01","00","00","00","00","00","01","00","01","00","01","00","01","00","01","00","00","00","00","00","01","00","01","00","01",
"00","01","00","01","00","01","00","00","00","00","00","01","00","01","00","01","00","01","00","01","00","00","00","00","00","01","00","01","00","00","00","00",
"00","01","01","01","01","00","01","00","01","00","00","00","01","00","01","00","01","00","01","00","01","00","01","00","00","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","00","00","01","00","01","00","01","00","01","00","01","00","01","00","00","00","01","00","01","00","00","00","00","00",
"00","01","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","00","00","00","00",
"00","01","01","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","00","00","00","00","00",
"00","01","01","00","00","01","01","01","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","00","00","00","01","01","00","00","00",
"00","01","00","00","00","00","01","01","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","00","00","01","01","01","01","00","00",
"00","01","00","00","00","00","01","01","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","00","00","01","01","01","01","00","00",
"00","01","01","00","00","01","01","01","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","00","00","00","01","01","00","00","00",
"00","01","01","01","01","01","01","01","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","01","01","00","00","01","01","01","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","01","01","00","00","00",
"00","01","00","00","00","00","01","01","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","01","01","01","01","00","00",
"00","01","00","00","00","00","01","01","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","01","01","01","01","00","00",
"00","01","01","00","00","01","01","01","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","01","01","00","00","00",
"00","01","01","01","01","01","01","01","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11",
"11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11",
"11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11",
"11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11",
"11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11",
"11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11",
"11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11",
"11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11",
"11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11",
"11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11",
"11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11",
"11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","00","00","00","00","00","00","00","00",
"00","01","01","00","00","01","01","01","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","00","00","00","01","01","00","00","00",
"00","01","00","00","00","00","01","01","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","00","00","01","01","01","01","00","00",
"00","01","00","00","00","00","01","01","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","00","00","01","01","01","01","00","00",
"00","01","01","00","00","01","01","01","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","00","00","00","01","01","00","00","00",
"00","01","01","01","01","01","01","01","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","01","01","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","01","01","00","00","01","01","01","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","01","01","00","00","00",
"00","01","00","00","00","00","01","01","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","01","01","01","01","00","00",
"00","01","00","00","00","00","01","01","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","01","01","01","01","00","00",
"00","01","01","00","00","01","01","01","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","01","01","00","00","00",
"00","01","01","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","01","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","01","01","01","01","00","00","00","00","01","01","00","00","00","00","00","00","00","00","00","00","00","00","01","01","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","01","01","00","00","00","00","00","00","00","00","00","00","00","00","01","01","00","00","00","00","00","00","00","00","00",
"00","01","01","01","00","00","00","00","01","01","01","01","00","00","00","00","00","00","00","00","00","00","01","01","01","01","00","00","00","00","00","00",
"00","00","00","00","00","00","01","01","01","01","00","00","00","00","00","00","00","00","00","00","01","01","01","01","00","00","00","00","00","00","00","00",
"00","01","01","00","00","00","00","00","01","01","01","01","00","00","00","00","00","00","00","00","00","00","01","01","01","01","00","00","00","00","00","00",
"00","00","00","00","00","00","01","01","01","01","00","00","00","00","00","00","00","00","00","00","01","01","01","01","00","00","00","00","00","00","00","00",
"00","01","00","00","00","00","00","00","00","01","01","00","00","00","00","00","00","00","00","00","00","00","00","01","01","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","01","01","00","00","00","00","00","00","00","00","00","00","00","00","01","01","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
-----------------------------------------------KONEC KAMENU/ZACATEK HRACE-------------------------------------
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00",
"00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11",
"11","11","11","11","11","00","00","10","10","10","10","10","10","10","10","00","00","00","00","11","11","11","11","11","11","11","11","11","00","00","00","00",
"00","00","00","11","11","11","11","11","11","11","11","11","11","11","00","00","00","01","00","00","00","00","00","11","11","11","11","11","11","11","11","11",
"11","11","11","11","00","00","10","10","10","10","10","10","10","10","10","10","10","10","00","00","11","11","11","11","11","11","11","11","11","00","00","00",
"00","00","00","11","11","11","11","11","11","11","11","11","11","00","01","00","00","00","00","00","00","01","00","00","00","11","11","11","11","11","11","11",
"11","11","11","11","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","11","11","11","11","11","11","11","00","00","00",
"00","00","11","11","11","11","11","11","11","11","11","11","00","00","00","10","10","10","10","10","10","00","00","00","00","00","00","11","11","11","11","11",
"11","11","11","00","00","00","10","10","10","10","10","10","10","00","00","10","10","10","10","10","10","10","00","00","11","11","11","11","11","11","00","00",
"00","00","11","11","11","11","11","11","11","11","11","00","00","00","10","10","10","10","10","10","10","10","10","00","01","00","00","11","11","11","11","11",
"11","11","11","00","00","10","00","10","10","10","10","10","10","00","00","00","00","10","10","10","10","10","10","10","00","00","11","11","11","11","00","00",
"00","00","11","11","11","11","11","11","11","11","00","00","00","10","10","10","10","01","01","01","01","10","10","10","00","00","00","11","11","11","11","11",
"11","11","00","00","10","10","00","10","10","10","10","10","10","00","00","00","00","00","00","10","10","10","10","10","10","10","00","11","11","11","00","00",
"00","00","11","11","11","11","11","11","11","00","01","00","10","10","10","01","01","01","01","01","01","01","10","10","10","00","00","00","11","11","11","11",
"11","11","00","00","10","10","00","00","10","10","10","10","10","10","00","00","00","00","00","00","00","10","10","10","10","10","10","00","11","11","00","00",
"00","11","11","11","11","11","11","11","11","00","00","00","10","10","01","01","01","01","10","10","10","10","10","10","10","00","01","00","11","11","11","11",
"11","11","00","00","10","00","00","00","00","10","10","10","10","10","10","00","00","00","00","00","00","00","10","10","10","10","10","00","11","11","11","00",
"00","11","11","11","11","11","11","11","11","00","00","10","10","01","01","01","01","10","10","10","10","10","10","10","10","10","00","00","11","11","11","11",
"11","11","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","00","00","00","00","00","00","10","10","10","10","10","00","11","11","00",
"00","11","11","11","11","11","11","11","11","00","00","10","01","01","01","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","11","11",
"11","11","00","00","00","00","00","00","00","10","00","00","00","10","10","10","10","10","10","10","00","00","00","10","10","10","10","10","00","11","11","00",
"00","11","11","11","11","11","11","11","00","01","00","10","01","01","10","10","10","10","10","10","10","10","10","10","10","10","10","00","01","00","11","11",
"11","11","11","00","00","00","00","00","10","10","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","11","00",
"00","11","11","11","11","11","11","11","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","11",
"11","11","11","00","00","00","00","00","10","00","00","00","00","00","10","00","00","00","10","10","10","10","10","10","10","10","10","10","10","00","11","00",
"00","11","11","11","11","11","11","11","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","11",
"11","11","11","11","00","00","00","00","00","00","00","00","00","00","10","10","00","00","00","00","10","10","10","10","10","10","10","10","00","11","11","00",
"00","11","11","11","11","11","11","11","00","00","10","10","01","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","11",
"11","11","11","11","11","00","00","00","00","00","00","00","00","10","10","00","00","00","00","00","00","00","00","10","10","10","00","00","00","11","11","00",
"00","11","11","11","11","11","11","00","00","00","10","01","01","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","01","00","11","11",
"11","11","11","11","11","11","00","00","00","00","00","00","00","10","10","00","00","00","00","00","10","10","10","00","00","00","00","00","00","11","11","00",
"00","11","11","11","11","11","11","00","01","00","10","01","01","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","11","11",
"11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","10","10","10","00","00","00","10","00","00","11","11","11","00",
"00","11","11","11","11","11","11","00","00","10","10","01","01","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","11","11","11","11",
"11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","10","10","00","00","00","00","10","00","00","11","11","11","00",
"00","11","11","11","11","11","11","00","00","10","10","01","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","11","11","11",
"11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","10","00","00","11","11","11","11","00",
"00","11","11","11","11","11","11","00","00","10","10","01","10","10","10","10","10","10","10","10","10","10","10","10","00","01","00","11","11","11","11","11",
"11","11","11","00","00","00","00","00","00","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","00",
"00","11","11","11","11","11","11","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","11","11","11","11",
"00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","00","00","00","00","00","00","00","00","11","11","11","11","11","11","00",
"00","11","11","11","11","11","11","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","11","11","11","11","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","00","00","00","11","11","11","11","11","11","11","11","00",
"00","11","11","11","11","11","11","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","00","01","00","11","11","11","11","11","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00",
"00","11","11","11","11","11","11","00","01","00","10","10","10","10","10","10","10","10","10","10","00","00","00","00","00","11","11","11","11","00","00","00",
"00","00","00","01","00","01","00","01","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00",
"00","11","11","11","11","11","11","11","00","00","10","10","10","10","10","10","10","10","00","00","00","00","00","11","11","11","11","11","00","00","00","00",
"00","00","01","00","01","00","01","00","01","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00",
"00","11","11","11","11","11","11","11","00","00","00","10","10","10","10","00","00","00","00","00","00","11","11","11","11","11","11","11","00","00","00","00",
"00","01","00","01","00","01","00","01","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00",
"00","11","11","11","11","11","11","11","11","00","00","00","00","00","00","01","00","00","00","11","11","11","11","11","11","11","11","00","00","00","00","00",
"01","00","01","00","01","00","01","00","00","00","00","00","01","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00",
"00","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","01",
"00","01","00","01","00","01","00","00","00","00","00","01","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00",
"00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","01","00",
"01","00","01","00","00","00","00","00","00","00","01","00","01","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","00",
"00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00",
"00","00","00","00","00","11","11","00","00","01","00","01","00","01","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","00",
"00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00",
"00","00","00","00","00","11","11","00","01","00","01","00","01","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","00",
"00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","01","00",
"01","00","01","00","00","00","00","00","00","01","00","01","00","01","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","00",
"00","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","01",
"00","01","00","01","00","01","00","00","00","00","01","00","01","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00",
"00","11","11","11","11","11","11","11","11","00","00","00","00","00","00","01","00","00","00","11","11","11","11","11","11","11","11","00","00","00","00","00",
"01","00","01","00","01","00","01","00","00","00","00","01","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00",
"00","11","11","11","11","11","11","11","00","00","00","10","10","10","10","00","00","00","00","00","00","11","11","11","11","11","11","00","00","00","00","00",
"00","01","00","01","00","01","00","01","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00",
"00","11","11","11","11","11","11","11","00","00","10","10","10","10","10","10","10","10","00","00","00","00","00","11","11","11","11","11","00","00","00","00",
"00","00","01","00","01","00","01","00","01","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00",
"00","11","11","11","11","11","11","00","01","00","10","01","01","01","01","01","01","10","10","10","00","00","00","00","00","11","11","11","11","00","00","00",
"00","00","00","01","00","01","00","01","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00",
"00","11","11","11","11","11","11","00","00","10","01","01","01","01","01","01","01","01","01","10","10","10","00","01","00","11","11","11","11","11","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00",
"00","11","11","11","11","11","11","00","00","10","01","01","10","10","10","10","10","10","01","01","01","10","10","00","00","00","11","11","11","11","11","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","00","00","00","11","11","11","11","11","11","11","11","00",
"00","11","11","11","11","11","11","00","00","10","10","10","10","10","10","10","10","10","10","01","01","01","10","10","00","00","00","11","11","11","11","11",
"00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","00","00","00","00","00","00","00","00","11","11","11","11","11","11","00",
"00","11","11","11","11","11","11","00","00","10","10","10","10","10","10","10","10","10","10","10","01","01","01","10","00","01","00","11","11","11","11","11",
"11","11","11","00","00","00","00","00","00","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","00",
"00","11","11","11","11","11","11","00","00","10","10","01","10","10","10","10","10","10","10","10","10","01","01","01","10","00","00","00","11","11","11","11",
"11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","10","00","00","11","11","11","11","00",
"00","11","11","11","11","11","11","00","00","10","10","01","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","11","11","11","11",
"11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","10","10","00","00","00","00","10","00","00","11","11","11","00",
"00","11","11","11","11","11","11","00","01","00","10","01","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","11","11",
"11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","10","10","10","00","00","00","10","00","00","11","11","11","00",
"00","11","11","11","11","11","11","00","00","00","10","01","01","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","01","00","11","11",
"11","11","11","11","11","11","00","00","00","00","00","00","00","10","10","00","00","00","00","00","10","10","10","00","00","00","00","00","00","11","11","00",
"00","11","11","11","11","11","11","11","00","00","10","01","01","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","11",
"11","11","11","11","11","00","00","00","00","00","00","00","00","10","10","00","00","00","00","00","00","00","00","10","10","10","00","00","00","11","11","00",
"00","11","11","11","11","11","11","11","00","00","10","10","01","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","11",
"11","11","11","11","00","00","00","00","00","00","00","00","00","00","10","10","00","00","00","00","10","10","10","10","10","10","10","10","00","11","11","00",
"00","11","11","11","11","11","11","11","00","00","10","10","01","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","11",
"11","11","11","00","00","00","00","00","10","00","00","00","00","00","10","00","00","00","10","10","10","10","10","10","10","10","10","10","10","00","11","00",
"00","11","11","11","11","11","11","11","00","01","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","01","00","11","11",
"11","11","11","00","00","00","00","00","10","10","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","11","00",
"00","11","11","11","11","11","11","11","11","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","11","11",
"11","11","00","00","00","00","00","00","00","10","00","00","00","10","10","10","10","10","10","10","00","00","00","10","10","10","10","10","00","11","11","00",
"00","11","11","11","11","11","11","11","11","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","11","11","11","11",
"11","11","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","00","00","00","00","00","00","10","10","10","10","10","00","11","11","00",
"00","11","11","11","11","11","11","11","11","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","00","01","00","11","11","11","11",
"11","11","00","00","10","00","00","00","00","10","10","10","10","10","10","00","00","00","00","00","00","00","10","10","10","10","10","00","11","11","11","00",
"00","00","11","11","11","11","11","11","11","00","01","00","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","11","11","11",
"11","11","00","00","10","10","00","00","10","10","10","10","10","10","00","00","00","00","00","00","00","10","10","10","10","10","10","00","11","11","00","00",
"00","00","11","11","11","11","11","11","11","11","00","00","00","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","11","11","11","11",
"11","11","00","00","10","10","00","10","10","10","10","10","10","00","00","00","00","00","00","10","10","10","10","10","10","10","00","11","11","11","00","00",
"00","00","11","11","11","11","11","11","11","11","11","00","00","00","10","10","10","10","10","10","10","10","10","00","01","00","00","11","11","11","11","11",
"11","11","11","00","00","10","00","10","10","10","10","10","10","00","00","00","00","10","10","10","10","10","10","10","00","00","11","11","11","11","00","00",
"00","00","11","11","11","11","11","11","11","11","11","11","00","00","00","10","10","10","10","10","10","00","00","00","00","00","00","11","11","11","11","11",
"11","11","11","00","00","00","10","10","10","10","10","10","10","00","00","10","10","10","10","10","10","10","00","00","11","11","11","11","11","11","00","00",
"00","00","00","11","11","11","11","11","11","11","11","11","11","00","01","00","00","00","00","00","00","01","00","00","00","11","11","11","11","11","11","11",
"11","11","11","11","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","11","11","11","11","11","11","11","00","00","00",
"00","00","00","11","11","11","11","11","11","11","11","11","11","11","00","00","00","01","00","00","00","00","00","11","11","11","11","11","11","11","11","11",
"11","11","11","11","00","00","10","10","10","10","10","10","10","10","10","10","10","10","00","00","11","11","11","11","11","11","11","11","11","00","00","00",
"00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11",
"11","11","11","11","11","00","00","10","10","10","10","10","10","10","10","00","00","00","00","11","11","11","11","11","11","11","11","11","00","00","00","00",
"00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
---------------------------------------------KONEC HRACE/ZACATEK JIDLA-----------------------------------------
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "01", "01", "01", "10", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", 
"11", "11", "11", "11", "11", "11", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", 
"11", "11", "11", "11", "11", "11", "11", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "10", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "11", "11", "11", "11", "11", 
"11", "11", "11", "11", "11", "11", "11", "11", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "10", "11", "10", "11", "11", 
"11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "10", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "11", "11", "11", "11", "11", 
"11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "10", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "11", "11", "11", "11", "11", "11", 
"11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "10", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "10", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "11", "11", "11", "11", "11", 
"11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "10", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "10", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "11", "11", "11", "11", "11", 
"11", "11", "11", "00", "00", "00", "11", "11", "11", "11", "11", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "10", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "11", "11", "11", "11", "11", 
"11", "11", "00", "00", "00", "00", "00", "00", "11", "11", "11", "11", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "10", "10", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "11", "11", "11", "11", "11", 
"11", "11", "00", "00", "00", "00", "00", "00", "00", "11", "11", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "10", "11", "10", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "11", "11", "11", "11", "11", 
"11", "11", "00", "00", "00", "00", "00", "00", "00", "00", "11", "11", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "10", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "10", "10", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "00", "00", "11", "11", "11", 
"11", "11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "10", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "10", "11", "10", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "00", "00", "00", "00", "11", "11", 
"11", "11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "10", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "10", "10", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "00", "00", "00", "00", "00", "11", 
"11", "11", "11", "11", "11", "00", "00", "00", "00", "00", "00", "00", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "10", "11", "10", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "11", "00", "00", "00", "00", "00", "00", "00", 
"11", "11", "00", "00", "00", "11", "00", "00", "00", "00", "00", "11", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "10", "10", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "00", "00", "00", "00", "00", "00", "00", 
"11", "00", "00", "00", "00", "00", "11", "11", "11", "11", "11", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "10", "11", "10", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "11", "00", "00", "00", "00", "00", "00", "00", 
"11", "00", "00", "00", "00", "00", "11", "11", "11", "11", "11", "11", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "10", "10", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "00", "00", "00", "00", "00", "00", "00", 
"11", "00", "00", "00", "00", "00", "11", "11", "11", "11", "11", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "10", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "10", "11", "10", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "11", "00", "00", "00", "00", "00", "00", "00", 
"11", "00", "00", "00", "00", "00", "11", "11", "11", "11", "11", "11", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "10", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "10", "10", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "00", "00", "00", "00", "00", "00", "00", 
"11", "11", "00", "00", "00", "11", "00", "00", "00", "00", "00", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "10", "11", "10", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "00", "00", "00", "00", "00", "11", 
"11", "11", "11", "11", "11", "00", "00", "00", "00", "00", "00", "00", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "10", "10", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "00", "00", "00", "00", "11", "11", 
"11", "11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "10", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "10", "11", "10", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "00", "00", "11", "11", "11", 
"11", "11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "10", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "10", "10", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "11", "11", "11", "11", "11", 
"11", "11", "00", "00", "00", "00", "00", "00", "00", "00", "11", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "10", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "10", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "11", "11", "11", "11", "11", 
"11", "11", "00", "00", "00", "00", "00", "00", "00", "11", "11", "11", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "01", "10", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "10", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "11", "11", "11", "11", "11", 
"11", "11", "00", "00", "00", "00", "00", "00", "11", "11", "11", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "01", "10", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "10", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "11", "11", "11", "11", "11", 
"11", "11", "11", "00", "00", "00", "11", "11", "11", "11", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "10", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "11", "11", "11", "11", 
"11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "10", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", 
"11", "10", "11", "11", "11", "11", "11", "11", "11", "11", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "10", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "11", "11", "11", "11", "11", 
"11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "10", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "11", "11", "11", "11", "11", 
"11", "11", "11", "11", "11", "11", "11", "11", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "10", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "11", "11", 
"11", "11", "11", "11", "11", "11", "11", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", 
"11", "11", "11", "11", "11", "11", "11", "10", "11", "10", "11", "10", "10", "10", "10", "10", "10", "10", "10", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "10", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", 
"00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
-------------------------------------------------------KONEC JIDLA/ZACATEK LOGA----------------------------------------------------------
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","10","10","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","10","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","10","10","00","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","10","00","00","10","10","10","10","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","11","11","11","11","11","11","11","11","11",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","11","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","11","11","01","01","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","11","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","11","11","01","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","11",
"00","00","00","00","00","00","00","00","00","00","00","00","11","11","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11",
"11","11","11","11","00","00","00","00","00","00","00","00","00","11","11","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","00","11","11","11","11","00","00","00","00","00","00","00","11","11","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11",
"11","11","11","11","00","00","00","00","00","00","00","00","00","11","11","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","11",
"00","00","00","00","00","00","00","00","00","00","00","00","11","11","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","11","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","11","11","01","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","11","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","11","11","01","01","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","11","11","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","11","11","11","11","11","11","11","11","11","11","11","11","11",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","00","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","11","11","11","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"00","00","00","00","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","11","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","00","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","00","11","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","00","11","00","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","00","11","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","00","11","00","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","11","11","11","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11",
"00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","10",
"00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11",
"00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","11",
"00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","11","00","00","00","00","00","00","00","00","00",
"00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","00","00","00","00","00","00",
"00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","11","00","00","00","00","00","00","00","00","00",
"00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","11",
"00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11",
"00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","10",
"11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11",
"11","00","11","00","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","00","11","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","00","11","00","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","00","11","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","00","11","00","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","00","11","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","00","11","00","11","11","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00",
"10","00","10","00","10","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11",
"11","11","11","11","11","11","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00",
"10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00",
"10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00",
"10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00",
"10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00",
"10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00",
"10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00",
"10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00",
"10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00",
"10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00",
"10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00",
"10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00",
"10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10",
"00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00",
"10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","10","10","00",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","10","10","10","10","10","10","10",
"10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","10","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","10","10","10","10","10","10","10",
"10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","10","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","10","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","10","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","10","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","10","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","10","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","10","00","00","00","00","00","00","00","00","00",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","10","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","10","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00",
"11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","00","10","00","10","00","10","00",
"10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","10","00","10","00","10","00","10",
"00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","11","11","11","11","11","11","00","11","00","11","00","11","00","11","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","11","11","11","11","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","11","11","11","11","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","11","11","11","11","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11",
"11","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","11","11","00","11",
"00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","11","11","00","00","00","00","00","11","00",
"11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","00","00","00","00","00","00","00","00","00","11","00","11",
"00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","11","11","11","11","11","00","11","00","11","00","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","11","00","11","00",
"11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","11","11","11","11","11","00","00","00","11","00","11","00","11","00","11","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","00","11","00","11","00","11",
"00","11","00","11","00","11","00","11","00","11","11","11","11","11","11","11","00","00","00","00","00","00","00","00","11","11","00","11","00","11","00","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","11","00","11","00","11","00",
"11","00","11","00","11","11","11","11","11","11","00","01","01","01","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","11","00","00","00","00","00","00","00","11","00","11","00","11","00","11",
"11","11","11","11","11","00","00","00","00","00","00","01","01","01","01","00","00","00","00","00","00","00","00","00","11","11","00","11","00","11","00","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","11","00","00","00","00","00","00","11","11","11","11","11","11","11","11",
"10","10","10","10","00","00","00","00","00","00","00","00","01","01","01","01","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","11","00","00","00","00","00","11","11","11","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","00","00","01","01","01","01","00","00","00","00","00","00","00","11","11","00","11","00","11","00","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","11","00","00","00","00","11","11","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","00","00","00","01","01","01","01","00","00","00","00","00","00","11","00","11","00","11","00","11","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","11","00","00","00","11","00","11","00","00","00","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","00","00","00","00","01","01","01","01","00","00","00","00","00","11","11","00","11","00","11","00","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","00","00","11","00","11","11","00","00","00","00","00","00","00","00",
"00","00","10","10","10","00","00","00","00","00","00","00","00","00","00","00","01","01","01","01","00","00","00","00","11","00","11","00","11","00","11","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","00","11","00","11","00","11","11","11","11","11","11","11","11","11",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","11","00","11","00","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","11","00","11","00","11","00","11","11","11","11","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","00","11","00","11","00","11","00","11","00","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","00","11","00","11","00","11","00","11","00","11","11","11","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","11",
"11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","00","11","00","11","00","11","00","11","00","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"00","11","00","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","00","11","00","11","00","11","00","11","00","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"11","00","11","00","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"00","11","00","11","00","11","00","11","11","11","00","00","00","00","00","00","00","00","00","01","11","11","00","11","00","11","00","11","00","11","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"11","00","11","00","11","00","11","00","11","11","11","11","00","00","00","00","00","00","01","01","11","11","11","11","11","11","11","11","11","11","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"00","11","00","11","00","11","00","11","00","11","00","11","11","11","00","00","00","01","01","01","01","00","00","00","00","00","00","00","00","11","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"11","00","11","00","11","00","11","00","11","00","11","00","11","11","11","11","01","01","01","01","00","00","00","00","00","00","00","00","00","11","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","11","00","11","00","11","00","11","00","11","11","11","11","11","11","11",
"00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","11","01","00","00","00","00","00","00","00","00","00","00","11","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","11","11","00","11","00","11","00","11","11","10","10","10","10","11","11",
"11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","11","11","00","00","00","00","00","00","00","00","00","11","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00","11","00","11","00","11","00","11","00","11","10","10","10","10","10","10",
"11","11","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","11","11","00","00","00","00","00","00","11","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","11","11","00","11","00","11","00","11","11","10","10","10","10","10","10",
"10","10","11","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","11","00","00","00","00","11","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","11","00","11","00","11","00","11","00","11","10","10","10","10","10","10",
"10","10","10","10","11","11","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","11","11","00","00","11","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","00","11","00","11","00","11","11","10","10","10","10","10","10",
"10","10","10","10","00","00","11","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","00","00","00","00","11","11","11","11","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","11","00","11","00","11","00","11","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","11","11","11","11","00","11","00","11","00","11","00","11","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","00","11","00","11","00","11","11","11","11","11","11","11","11",
"11","11","11","10","00","00","00","00","00","00","00","11","11","11","11","00","11","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"00","11","11","10","00","00","00","00","00","00","00","01","01","11","11","11","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"11","00","11","10","00","00","00","00","00","00","00","01","01","01","00","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"00","11","11","10","00","00","00","00","00","00","00","01","01","01","00","00","00","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"11","00","11","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","11","11","11","11","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"00","11","11","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","11","11","11","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"11","00","11","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","11","11","11","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"00","11","11","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","01","00","11","11","11","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"11","11","11","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","01","00","00","00","11","11","11","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","11","11","11","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"11","00","11","00","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00","11",
"00","11","00","11","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00","11","00",
"11","00","11","00","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00","11","00","11",
"00","11","00","11","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00",
"11","00","11","00","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"00","11","00","11","00","11","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"11","00","11","00","11","11","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"11","11","11","11","11","11","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","11","00",
"11","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","00","00","00","00","00","00","11","10","10","10","10","00","00","00","00","00","10","10","10","10","10","11","00","11","00","11",
"11","00","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","00","11","00","00","00","00","00","00","00","11","00","00","00","00","00","00","00","00","10","10","10","10","10","10","11","11","00","11","00",
"11","00","00","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","00","00","11","00","00","00","00","00","00","00","11","00","00","00","00","00","00","00","00","10","10","10","10","10","10","11","00","11","00","11",
"11","00","00","00","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","00","00","00","11","00","00","00","00","00","00","00","11","00","00","00","00","00","00","00","00","10","10","10","10","10","10","11","11","00","11","00",
"11","01","00","00","00","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"00","00","00","00","11","00","00","00","00","00","00","11","11","00","00","00","00","00","00","00","00","10","10","10","10","10","10","11","00","11","00","11",
"11","01","01","00","00","00","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00",
"00","00","00","01","11","00","00","00","00","00","11","00","11","00","00","00","00","00","00","00","10","10","10","10","10","10","10","11","11","00","11","00",
"11","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00",
"00","00","01","01","11","00","00","00","00","11","00","11","11","00","00","00","00","00","00","00","10","10","10","10","10","10","10","11","00","11","00","11",
"11","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00",
"00","01","01","01","11","00","00","00","11","00","11","00","11","00","00","00","00","00","00","00","10","10","10","10","10","10","10","11","11","00","11","00",
"11","00","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","00","00","00","00",
"01","01","01","00","11","00","00","11","00","11","00","11","11","00","00","00","00","00","00","00","10","10","10","10","10","10","10","11","00","11","00","11",
"11","11","11","11","11","11","01","00","00","00","00","00","00","00","00","00","00","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","01","01","11","00","11","00","11","00","11","00","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","11","11","00","11","00",
"11","00","11","00","11","11","01","01","00","00","00","00","00","00","00","00","00","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","01","01","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","00","00","00","00","11","00","11","00","11",
"00","11","00","11","00","11","01","01","01","00","00","00","00","00","00","00","00","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","01","01","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","00","00","00","00","00","11","11","00","11","00",
"11","00","11","00","11","11","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"01","01","01","00","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","00","00","00","00","11","00","11","00","11",
"00","11","00","11","00","11","00","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","01","01","01","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","00","00","00","00","00","11","11","00","11","00",
"11","00","11","00","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","01","01","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","00","00","00","00","11","11","11","11","11",
"00","11","00","11","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","01","11","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","00","00","00","00","00","10","10","10","10","10",
"11","00","11","00","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","01","11","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","00","00","00","10","10","10","10","10","10",
"11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","01","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","10","10","10","10","10","10","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10",
"11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"00","11","00","11","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","11","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"11","00","11","00","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","11","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"00","11","00","00","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","01","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"11","00","00","00","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","01","01","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"00","00","00","00","00","11","00","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","01","01","01","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"00","00","00","00","00","11","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"01","01","01","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"00","00","00","00","00","11","01","01","01","00","00","00","00","00","00","00","00","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","01","01","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"00","00","00","00","00","11","01","01","00","00","00","00","00","00","00","00","00","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","01","01","11","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"00","00","00","00","00","11","01","00","00","00","00","00","00","00","00","00","00","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","01","01","01","01","11","11","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"00","00","00","00","00","11","00","00","00","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","00","00","00","00",
"01","01","01","00","00","00","00","00","00","11","11","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"00","00","00","00","00","11","00","00","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","00","00","00",
"00","01","01","01","00","00","00","00","00","00","00","00","11","11","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"00","00","00","00","00","11","00","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","00",
"00","00","01","01","01","00","00","00","00","00","00","00","00","00","00","11","11","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"00","00","00","00","00","11","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00",
"00","00","00","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","00","11","00","11","00","11","00","11","00","11",
"00","00","00","00","00","11","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"00","00","00","00","01","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","00","11","00","11","00","11","00",
"00","00","00","00","00","11","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","00","00","00","00","01","01","01","01","01","01","00","00","00","00","00","00","00","00","00","00","10","10","10","11","11","11","11","00","11","00","11",
"00","00","00","00","00","11","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","10","10","10","10","10","10","11","11","11","11","00",
"00","00","00","00","00","11","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","00","00","00","00","00","00","00","00","00","10","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","11","11",
"00","00","00","00","00","11","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"00","00","00","00","00","11","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"00","00","00","00","00","11","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"00","00","00","00","00","11","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"00","00","00","00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"00","00","00","00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"00","00","00","00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"00","00","00","00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","11","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"11","11","11","11","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","10","10","10","10","10","10","00","10","00",
"00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","11","10","10","10","10","10","10","00","10",
"00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","11","10","10","10","10","10","10","00",
"10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","10","10","10","10","10","00","10",
"00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","10","10","10","10","10","10","00",
"10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","10","10","10","10","10","10","10",
"00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","10","10","10","10","10","10","00",
"10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","10","10","10","10","10","10","10",
"00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","11","00","11","00","11","00","11","10","10","10","10","10","10","10",
"10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","00","11","00","11","00","11","11","10","10","10","10","10","10","10",
"10","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","11","00","11","00","11","00","11","10","10","10","10","10","10","10",
"10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","00","11","00","11","00","11","11","10","10","10","10","10","10","10",
"10","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","11","00","11","00","11","00","11","10","10","10","10","10","10","10",
"10","10","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","00","11","00","11","00","11","11","10","10","10","10","10","10","10",
"10","10","10","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","11","00","11","00","11","00","11","10","10","10","10","10","10","10",
"10","10","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","00","11","00","11","00","11","11","10","10","10","10","10","10","10",
"10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","11","00","11","00","11","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","00","11","00","11","00","11","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00",
"11","11","10","10","10","10","10","11","11","11","11","11","11","11","11","11","11","00","11","00","11","00","11","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00",
"00","11","10","10","10","10","10","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00",
"11","11","10","10","10","10","10","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00",
"00","11","10","10","10","10","10","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00",
"11","11","10","10","10","10","10","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00",
"11","11","10","10","10","10","10","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00",
"10","10","10","10","10","10","10","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00",
"10","10","10","10","10","10","10","11","00","11","00","11","00","11","00","11","00","00","00","11","00","11","11","11","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00",
"10","10","10","10","10","10","10","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00",
"00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00",
"11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00",
"00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00",
"11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00",
"00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00",
"11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00",
"00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00",
"11","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00",
"00","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00",
"11","00","11","11","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","00","11","00","11","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","00","11","00","11","00","11","11","11","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","00","11","00","11","00","11","00","11","11","11","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","00","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","00","11","00","11","00","11","00","11","00","11","00","00","11","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","00","11","00","11","00","11","00","11","00","00","00","00","00","11","11","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","00","11","00","11","00","11","00","11","00","00","00","00","00","00","00","00","00","11","11","11","11","10","10","10","10","10","10","10","10","10","10",
"10","10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","00","11","00","11","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","10","10","10","10","10","10","10","10",
"10","00","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","00","11","00","11","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","10","10","10","10","10","10","10",
"10","10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","00","11","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","00","11","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"00","10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","10","00",
"10","00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"00","10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","10","00",
"10","00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","00","10",
"00","10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","10","00",
"10","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","10","10","10","10","10","00","10",
"00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00",
"00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","00","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"11","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","00","11","00","11","00","11","00","11","00","11","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","00","00","00","00","00","00","00","00","11","11","11","11","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","00","00","00","00","00","00","11","11","11","00","00","11","11","11","11","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","00","00","00","11","11","11","11","00","00","00","00","00","00","00","11","11","11","11","00","00","01","01","01","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","01","01","01","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11",
"11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","11","11","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","11","11","11","11","01","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","11","11","11","11","00","00","01","01","01","00","00","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","11","11","11","00","00","00","00","00","01","01","01","00","00","00","00","11","11","11","11","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","11",
"11","11","11","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","11","11","11","11","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","11","11","11",
"10","10","00","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","11","11","11","11","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","11","11","11","11","10","10",
"10","10","00","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","01","00","00","11","11","11","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","11","11","11","11","10","10","10","10","10",
"10","10","00","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","11","11","11",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","11","11","11","11","10","10","10","10","10","10","10","10",
"10","10","00","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","11","11","11","10","10","10","10","10","10","10","10","10","10","10",
"10","10","00","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","00","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","10","00","00","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","10","10","00","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","01","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","01","10","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","01","10","10","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"11","11","11","11","11","11","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","11","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","00","00","00","00","00","00","00",
"00","00","00","00","00","11","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00",
"10","00","10","00","11","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","11","00","11","00","11","00","11","00","11","00","11","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","11","11","00","11","00","11","00","11","00","11","00","11","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","11","00","11","00","11","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00",
"11","11","11","11","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","11","11","00","11","00","11","00","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","00","00","00","00",
"00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","11","00","11","00","11","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00",
"00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","11","00","11","00","11","00","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00",
"00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","11","00","11","00","11","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00",
"00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","11","00","11","00","11","00","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00",
"00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","11","00","11","00","11","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00",
"00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","11","00","11","00","11","00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00",
"00","00","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","11","00","11","00","00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00",
"11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","11","00","11","00","00","00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00",
"00","11","11","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","11","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00",
"00","00","00","00","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","00","00","00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","11","11","11","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","11","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","10","11","11","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
"00","00","10","10","10","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","00","00","00","00","00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"11","11","00","10","00","10","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","00","10","00","10","00","10",
"00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","11","11","00","10","00","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","10","00","10","00","10","00",
"10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","00","00","00","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","00","00","00","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","10","10","10","10","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","00","00","00","00","00","00","00","00","00","00","00","00","00","11","00","00","00","00","00","00","00","11","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","10","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","10","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","10","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","10","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","10","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","10","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","10","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","10","10","10","10","10","10","10",
"10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","10","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","11","10","10","10","10","10","10","10","10",
"10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","10","00","00","00","00",
"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","10","10","10","10","10","10","10","10","10",
"10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","10","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","10","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","10","10","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00",
"10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10",
"00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00",
"10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00",
"10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00",
"10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00",
"10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00",
"10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00",
"10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00",
"10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00",
"10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","10","10","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00",
"10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00","00",
"10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00",
"10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00","00",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10",
"00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","10","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
---------------------------------------------------------KONEC LOGA/ZACATEK ENTERU-----------------------------------------------------
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"01","01","01","01","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","00","01","00","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","00","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00","01","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","01","00","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00","00",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
"01","01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"00","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","01","01","01","01","01","01","01","01",
"01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","01","01","00","01","01","00","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","01","01","00","01","01","00","01","01","01","01","01","01","00","00",
"00","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","01","01","01","01","01","00","01","01","01","01","01","00","00","00",
"00","00","00","01","01","01","01","01","01","01","01","01","01","00","00","01","01","00","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","01","01","01","01","01","00","01","01","01","01","00","00","00","00",
"00","00","00","00","01","01","01","01","01","01","01","01","00","01","01","00","01","01","00","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","00","01","01","00","01","01","00","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","00","01","01","00","01","01","00","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","01","00","01","01","00","00","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","00","00","01","01","01","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00","00","00","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","01","00","00","00","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","00","01","01","00","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","01","00","00","00","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","01","01","00","01","01","00","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00","00","00","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","01","01","00","01","01","00","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","01","01","01","01","01","00","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","01","01","01","01","01","00","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","00","01","01","00","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","00","01","01","00","00","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","00","01","01","00","01","00","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","01","01","00","01","01","01","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","01","00","00","01","01","01","00","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","01","01","00","00","01","01","01","01","01","01","01","01","01","00",
"00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","00","01","01","00","01","00","01","01","01","01","00","00","00","00","00",
"00","01","01","01","01","01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","00","00","01","01","01","00","01","01","01","00","00","00","00","00",
"00","01","01","01","01","01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","01","01","01","01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","01","01","01","01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","00","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","00","00","00","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01",
"01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"01","01","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"01","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
--------------------------------------------------KONEC ENTERU/ZACATEK SIPKY--------------------------------------------------
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", 
"01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00"
------------------------------------------------------------KONEC SIPKY------------------------------------------------
);

signal y_x1, y_x2 : std_logic_vector(15 downto 0) := (others => '0');

begin

	y_x1 <= address_y1 & address_x1;
	y_x2 <= address_y2 & address_x2;

	process (clock)
	begin
   if (rising_edge(clock)) then
      if (en = '1') then
         if (we = '1') then
            rom(to_integer(unsigned(y_x1))) <= data_in;
         end if;
          data_out1 <= rom(to_integer(unsigned(y_x1)));
			 data_out2 <= rom(to_integer(unsigned(y_x2)));
      end if;
   end if;
end process;


end Behavioral;

